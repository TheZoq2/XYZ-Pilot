library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Datatypes;

entity sin_table is
    port(
            angle: in unsigned(7 downto 0);
            result:  out datatypes.small_number_t
        );
end entity;

architecture behaviour of sin_table is
begin
    with angle select
        result <= x"0000" when x"00",
x"0003" when x"01",
x"0006" when x"02",
x"0009" when x"03",
x"000c" when x"04",
x"000f" when x"05",
x"0012" when x"06",
x"0016" when x"07",
x"0019" when x"08",
x"001c" when x"09",
x"001f" when x"0a",
x"0022" when x"0b",
x"0025" when x"0c",
x"0028" when x"0d",
x"002b" when x"0e",
x"002f" when x"0f",
x"0032" when x"10",
x"0035" when x"11",
x"0038" when x"12",
x"003b" when x"13",
x"003e" when x"14",
x"0041" when x"15",
x"0044" when x"16",
x"0047" when x"17",
x"004a" when x"18",
x"004d" when x"19",
x"0050" when x"1a",
x"0053" when x"1b",
x"0056" when x"1c",
x"0059" when x"1d",
x"005c" when x"1e",
x"005f" when x"1f",
x"0062" when x"20",
x"0065" when x"21",
x"0068" when x"22",
x"006a" when x"23",
x"006d" when x"24",
x"0070" when x"25",
x"0073" when x"26",
x"0076" when x"27",
x"0079" when x"28",
x"007b" when x"29",
x"007e" when x"2a",
x"0081" when x"2b",
x"0084" when x"2c",
x"0086" when x"2d",
x"0089" when x"2e",
x"008c" when x"2f",
x"008e" when x"30",
x"0091" when x"31",
x"0093" when x"32",
x"0096" when x"33",
x"0099" when x"34",
x"009b" when x"35",
x"009e" when x"36",
x"00a0" when x"37",
x"00a2" when x"38",
x"00a5" when x"39",
x"00a7" when x"3a",
x"00aa" when x"3b",
x"00ac" when x"3c",
x"00ae" when x"3d",
x"00b1" when x"3e",
x"00b3" when x"3f",
x"00b5" when x"40",
x"00b7" when x"41",
x"00b9" when x"42",
x"00bc" when x"43",
x"00be" when x"44",
x"00c0" when x"45",
x"00c2" when x"46",
x"00c4" when x"47",
x"00c6" when x"48",
x"00c8" when x"49",
x"00ca" when x"4a",
x"00cc" when x"4b",
x"00ce" when x"4c",
x"00d0" when x"4d",
x"00d1" when x"4e",
x"00d3" when x"4f",
x"00d5" when x"50",
x"00d7" when x"51",
x"00d8" when x"52",
x"00da" when x"53",
x"00dc" when x"54",
x"00dd" when x"55",
x"00df" when x"56",
x"00e0" when x"57",
x"00e2" when x"58",
x"00e3" when x"59",
x"00e5" when x"5a",
x"00e6" when x"5b",
x"00e7" when x"5c",
x"00e9" when x"5d",
x"00ea" when x"5e",
x"00eb" when x"5f",
x"00ec" when x"60",
x"00ee" when x"61",
x"00ef" when x"62",
x"00f0" when x"63",
x"00f1" when x"64",
x"00f2" when x"65",
x"00f3" when x"66",
x"00f4" when x"67",
x"00f5" when x"68",
x"00f6" when x"69",
x"00f7" when x"6a",
x"00f7" when x"6b",
x"00f8" when x"6c",
x"00f9" when x"6d",
x"00fa" when x"6e",
x"00fa" when x"6f",
x"00fb" when x"70",
x"00fb" when x"71",
x"00fc" when x"72",
x"00fc" when x"73",
x"00fd" when x"74",
x"00fd" when x"75",
x"00fe" when x"76",
x"00fe" when x"77",
x"00fe" when x"78",
x"00ff" when x"79",
x"00ff" when x"7a",
x"00ff" when x"7b",
x"00ff" when x"7c",
x"00ff" when x"7d",
x"00ff" when x"7e",
x"00ff" when x"7f",
x"00ff" when x"80",
x"00ff" when x"81",
x"00ff" when x"82",
x"00ff" when x"83",
x"00ff" when x"84",
x"00ff" when x"85",
x"00ff" when x"86",
x"00fe" when x"87",
x"00fe" when x"88",
x"00fe" when x"89",
x"00fd" when x"8a",
x"00fd" when x"8b",
x"00fc" when x"8c",
x"00fc" when x"8d",
x"00fb" when x"8e",
x"00fb" when x"8f",
x"00fa" when x"90",
x"00fa" when x"91",
x"00f9" when x"92",
x"00f8" when x"93",
x"00f7" when x"94",
x"00f7" when x"95",
x"00f6" when x"96",
x"00f5" when x"97",
x"00f4" when x"98",
x"00f3" when x"99",
x"00f2" when x"9a",
x"00f1" when x"9b",
x"00f0" when x"9c",
x"00ef" when x"9d",
x"00ee" when x"9e",
x"00ec" when x"9f",
x"00eb" when x"a0",
x"00ea" when x"a1",
x"00e9" when x"a2",
x"00e7" when x"a3",
x"00e6" when x"a4",
x"00e5" when x"a5",
x"00e3" when x"a6",
x"00e2" when x"a7",
x"00e0" when x"a8",
x"00df" when x"a9",
x"00dd" when x"aa",
x"00dc" when x"ab",
x"00da" when x"ac",
x"00d8" when x"ad",
x"00d7" when x"ae",
x"00d5" when x"af",
x"00d3" when x"b0",
x"00d1" when x"b1",
x"00d0" when x"b2",
x"00ce" when x"b3",
x"00cc" when x"b4",
x"00ca" when x"b5",
x"00c8" when x"b6",
x"00c6" when x"b7",
x"00c4" when x"b8",
x"00c2" when x"b9",
x"00c0" when x"ba",
x"00be" when x"bb",
x"00bc" when x"bc",
x"00b9" when x"bd",
x"00b7" when x"be",
x"00b5" when x"bf",
x"00b3" when x"c0",
x"00b1" when x"c1",
x"00ae" when x"c2",
x"00ac" when x"c3",
x"00aa" when x"c4",
x"00a7" when x"c5",
x"00a5" when x"c6",
x"00a2" when x"c7",
x"00a0" when x"c8",
x"009e" when x"c9",
x"009b" when x"ca",
x"0099" when x"cb",
x"0096" when x"cc",
x"0093" when x"cd",
x"0091" when x"ce",
x"008e" when x"cf",
x"008c" when x"d0",
x"0089" when x"d1",
x"0086" when x"d2",
x"0084" when x"d3",
x"0081" when x"d4",
x"007e" when x"d5",
x"007b" when x"d6",
x"0079" when x"d7",
x"0076" when x"d8",
x"0073" when x"d9",
x"0070" when x"da",
x"006d" when x"db",
x"006a" when x"dc",
x"0068" when x"dd",
x"0065" when x"de",
x"0062" when x"df",
x"005f" when x"e0",
x"005c" when x"e1",
x"0059" when x"e2",
x"0056" when x"e3",
x"0053" when x"e4",
x"0050" when x"e5",
x"004d" when x"e6",
x"004a" when x"e7",
x"0047" when x"e8",
x"0044" when x"e9",
x"0041" when x"ea",
x"003e" when x"eb",
x"003b" when x"ec",
x"0038" when x"ed",
x"0035" when x"ee",
x"0032" when x"ef",
x"002f" when x"f0",
x"002b" when x"f1",
x"0028" when x"f2",
x"0025" when x"f3",
x"0022" when x"f4",
x"001f" when x"f5",
x"001c" when x"f6",
x"0019" when x"f7",
x"0016" when x"f8",
x"0012" when x"f9",
x"000f" when x"fa",
x"000c" when x"fb",
x"0009" when x"fc",
x"0006" when x"fd",
x"0003" when x"fe",
        x"0000" when others;
end architecture;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Datatypes;

entity cos_table is
    port(
            angle: in unsigned(7 downto 0);
            result:  out datatypes.small_number_t
        );
end entity;

architecture behaviour of cos_table is
begin
    with angle select
        result <= x"0100" when x"00",
        x"00ff" when x"01",
        x"00ff" when x"02",
        x"00ff" when x"03",
        x"00ff" when x"04",
        x"00ff" when x"05",
        x"00ff" when x"06",
        x"00ff" when x"07",
        x"00fe" when x"08",
        x"00fe" when x"09",
        x"00fe" when x"0a",
        x"00fd" when x"0b",
        x"00fd" when x"0c",
        x"00fc" when x"0d",
        x"00fc" when x"0e",
        x"00fb" when x"0f",
        x"00fb" when x"10",
        x"00fa" when x"11",
        x"00f9" when x"12",
        x"00f9" when x"13",
        x"00f8" when x"14",
        x"00f7" when x"15",
        x"00f6" when x"16",
        x"00f5" when x"17",
        x"00f4" when x"18",
        x"00f3" when x"19",
        x"00f2" when x"1a",
        x"00f1" when x"1b",
        x"00f0" when x"1c",
        x"00ef" when x"1d",
        x"00ee" when x"1e",
        x"00ed" when x"1f",
        x"00ec" when x"20",
        x"00eb" when x"21",
        x"00e9" when x"22",
        x"00e8" when x"23",
        x"00e7" when x"24",
        x"00e5" when x"25",
        x"00e4" when x"26",
        x"00e3" when x"27",
        x"00e1" when x"28",
        x"00e0" when x"29",
        x"00de" when x"2a",
        x"00dc" when x"2b",
        x"00db" when x"2c",
        x"00d9" when x"2d",
        x"00d7" when x"2e",
        x"00d6" when x"2f",
        x"00d4" when x"30",
        x"00d2" when x"31",
        x"00d0" when x"32",
        x"00cf" when x"33",
        x"00cd" when x"34",
        x"00cb" when x"35",
        x"00c9" when x"36",
        x"00c7" when x"37",
        x"00c5" when x"38",
        x"00c3" when x"39",
        x"00c1" when x"3a",
        x"00bf" when x"3b",
        x"00bd" when x"3c",
        x"00bb" when x"3d",
        x"00b8" when x"3e",
        x"00b6" when x"3f",
        x"00b4" when x"40",
        x"00b2" when x"41",
        x"00af" when x"42",
        x"00ad" when x"43",
        x"00ab" when x"44",
        x"00a8" when x"45",
        x"00a6" when x"46",
        x"00a4" when x"47",
        x"00a1" when x"48",
        x"009f" when x"49",
        x"009c" when x"4a",
        x"009a" when x"4b",
        x"0097" when x"4c",
        x"0095" when x"4d",
        x"0092" when x"4e",
        x"0090" when x"4f",
        x"008d" when x"50",
        x"008a" when x"51",
        x"0088" when x"52",
        x"0085" when x"53",
        x"0082" when x"54",
        x"0080" when x"55",
        x"007d" when x"56",
        x"007a" when x"57",
        x"0077" when x"58",
        x"0074" when x"59",
        x"0072" when x"5a",
        x"006f" when x"5b",
        x"006c" when x"5c",
        x"0069" when x"5d",
        x"0066" when x"5e",
        x"0063" when x"5f",
        x"0060" when x"60",
        x"005d" when x"61",
        x"005b" when x"62",
        x"0058" when x"63",
        x"0055" when x"64",
        x"0052" when x"65",
        x"004f" when x"66",
        x"004c" when x"67",
        x"0049" when x"68",
        x"0046" when x"69",
        x"0043" when x"6a",
        x"003f" when x"6b",
        x"003c" when x"6c",
        x"0039" when x"6d",
        x"0036" when x"6e",
        x"0033" when x"6f",
        x"0030" when x"70",
        x"002d" when x"71",
        x"002a" when x"72",
        x"0027" when x"73",
        x"0024" when x"74",
        x"0021" when x"75",
        x"001d" when x"76",
        x"001a" when x"77",
        x"0017" when x"78",
        x"0014" when x"79",
        x"0011" when x"7a",
        x"000e" when x"7b",
        x"000b" when x"7c",
        x"0007" when x"7d",
        x"0004" when x"7e",
        x"0001" when x"7f",
        x"8001" when x"80",
        x"8004" when x"81",
        x"8007" when x"82",
        x"800b" when x"83",
        x"800e" when x"84",
        x"8011" when x"85",
        x"8014" when x"86",
        x"8017" when x"87",
        x"801a" when x"88",
        x"801d" when x"89",
        x"8021" when x"8a",
        x"8024" when x"8b",
        x"8027" when x"8c",
        x"802a" when x"8d",
        x"802d" when x"8e",
        x"8030" when x"8f",
        x"8033" when x"90",
        x"8036" when x"91",
        x"8039" when x"92",
        x"803c" when x"93",
        x"803f" when x"94",
        x"8043" when x"95",
        x"8046" when x"96",
        x"8049" when x"97",
        x"804c" when x"98",
        x"804f" when x"99",
        x"8052" when x"9a",
        x"8055" when x"9b",
        x"8058" when x"9c",
        x"805b" when x"9d",
        x"805d" when x"9e",
        x"8060" when x"9f",
        x"8063" when x"a0",
        x"8066" when x"a1",
        x"8069" when x"a2",
        x"806c" when x"a3",
        x"806f" when x"a4",
        x"8072" when x"a5",
        x"8074" when x"a6",
        x"8077" when x"a7",
        x"807a" when x"a8",
        x"807d" when x"a9",
        x"807f" when x"aa",
        x"8082" when x"ab",
        x"8085" when x"ac",
        x"8088" when x"ad",
        x"808a" when x"ae",
        x"808d" when x"af",
        x"8090" when x"b0",
        x"8092" when x"b1",
        x"8095" when x"b2",
        x"8097" when x"b3",
        x"809a" when x"b4",
        x"809c" when x"b5",
        x"809f" when x"b6",
        x"80a1" when x"b7",
        x"80a4" when x"b8",
        x"80a6" when x"b9",
        x"80a8" when x"ba",
        x"80ab" when x"bb",
        x"80ad" when x"bc",
        x"80af" when x"bd",
        x"80b2" when x"be",
        x"80b4" when x"bf",
        x"80b6" when x"c0",
        x"80b8" when x"c1",
        x"80bb" when x"c2",
        x"80bd" when x"c3",
        x"80bf" when x"c4",
        x"80c1" when x"c5",
        x"80c3" when x"c6",
        x"80c5" when x"c7",
        x"80c7" when x"c8",
        x"80c9" when x"c9",
        x"80cb" when x"ca",
        x"80cd" when x"cb",
        x"80cf" when x"cc",
        x"80d0" when x"cd",
        x"80d2" when x"ce",
        x"80d4" when x"cf",
        x"80d6" when x"d0",
        x"80d7" when x"d1",
        x"80d9" when x"d2",
        x"80db" when x"d3",
        x"80dc" when x"d4",
        x"80de" when x"d5",
        x"80e0" when x"d6",
        x"80e1" when x"d7",
        x"80e3" when x"d8",
        x"80e4" when x"d9",
        x"80e5" when x"da",
        x"80e7" when x"db",
        x"80e8" when x"dc",
        x"80e9" when x"dd",
        x"80eb" when x"de",
        x"80ec" when x"df",
        x"80ed" when x"e0",
        x"80ee" when x"e1",
        x"80ef" when x"e2",
        x"80f0" when x"e3",
        x"80f1" when x"e4",
        x"80f2" when x"e5",
        x"80f3" when x"e6",
        x"80f4" when x"e7",
        x"80f5" when x"e8",
        x"80f6" when x"e9",
        x"80f7" when x"ea",
        x"80f8" when x"eb",
        x"80f9" when x"ec",
        x"80f9" when x"ed",
        x"80fa" when x"ee",
        x"80fb" when x"ef",
        x"80fb" when x"f0",
        x"80fc" when x"f1",
        x"80fc" when x"f2",
        x"80fd" when x"f3",
        x"80fd" when x"f4",
        x"80fe" when x"f5",
        x"80fe" when x"f6",
        x"80fe" when x"f7",
        x"80ff" when x"f8",
        x"80ff" when x"f9",
        x"80ff" when x"fa",
        x"80ff" when x"fb",
        x"80ff" when x"fc",
        x"80ff" when x"fd",
        x"80ff" when x"fe",
        x"8100" when others;
end architecture;
