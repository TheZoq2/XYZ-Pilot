
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Vector;

--Constants
package GPU_Info is
    --TODO: Optimse the size of obj addr and model addr
    --The length of the addresses and data in the object memory
    constant OBJ_ADDR_SIZE: positive := 9;
    constant OBJ_DATA_SIZE: positive := Vector.MEMORY_SIZE;

    subtype ObjAddr_t is unsigned(OBJ_ADDR_SIZE - 1 downto 0);
    subtype ObjData_t is std_logic_vector(OBJ_DATA_SIZE - 1 downto 0);

    constant MODEL_ADDR_SIZE: positive := 9;

    subtype ModelAddr_t is unsigned(MODEL_ADDR_SIZE - 1 downto 0);
    subtype ModelData_t is Vector.InMemory_t;
end package;

library IEEE;

use IEEE.Numeric_std.all;
use IEEE.std_logic_1164.all;

use work.Vector;
use work.GPU_Info;

entity ModelMem is
port (
        clk : in std_logic;
        -- port 1
        read_addr : in GPU_Info.ModelAddr_t;
        read_data : out GPU_Info.ModelData_t
    );
end entity;

architecture Behavioral of ModelMem is

-- Deklaration av ett dubbelportat block-RAM
-- med 2048 adresser av 8 bitars bredd.
type ram_t is array (0 to 511) of Vector.InMemory_t;

    -- Nollställ alla bitar på alla adresser
    signal ram : ram_t := ( 
    -- Start of ship
    0 => x"fff00000fffc0000",
    1 => x"fff0000000020000",
    2 => x"00170000ffff0000",
    3 => x"fff00000fffc0000",
    4 => x"0005fff8ffff0000",
    5 => x"00170000ffff0000",
    6 => x"0005000000010000",
    7 => x"00170000ffff0000",
    8 => x"fff00000fffc0000",
    9 => x"fff3fff3ffff0000",
    10 => x"fff3fff3ffff0000",
    11 => x"fff0000000020000",
    12 => x"fff3fff3ffff0000",
    13 => x"0005fff8ffff0000",
    14 => x"fff0000000020000",
    15 => x"fff8000000020000",
    16 => x"0001000000040000",
    17 => x"0005000000010000",
    18 => x"0005000000010000",
    19 => x"fffffffd00000000",
    20 => x"fff8000000020000",
    21 => x"fffcfffd00010000",
    22 => x"fffffffd00000000",
    23 => x"fffcfffd00010000",
    24 => x"fff8000000020000",
    25 => x"fffc000000040000",
    26 => x"fffc000000040000",
    27 => x"0001000000040000",
    28 => x"fffcfffd00010000",
    29 => x"fffc000000040000",
    30 => x"fffffffd00000000",
    31 => x"0001000000040000",
    32 => x"0005fff8ffff0000",
    33 => x"000cfff8ffff0000",
    34 => x"fff1fffdfffe0000",
    35 => x"fff1fffd00010000",
    36 => x"fff1fffdfffe0000",
    37 => x"fff2fff6ffff0000",
    38 => x"fff2fff6ffff0000",
    39 => x"fff1fffd00010000",
    40 => x"fff0000000020000",
    41 => x"fff1fffd00010000",
    42 => x"fff2fff6ffff0000",
    43 => x"fff3fff3ffff0000",
    44 => x"fff1fffdfffe0000",
    45 => x"fff00000fffc0000",
    46 => x"ffeefffcfffe0000",
    47 => x"ffeefffc00010000",
    48 => x"ffeefffcfffe0000",
    49 => x"ffeffff6ffff0000",
    50 => x"ffeffff6ffff0000",
    51 => x"ffeefffc00010000",
    52 => x"fff1fffd00010000",
    53 => x"ffeefffc00010000",
    54 => x"ffeffff6ffff0000",
    55 => x"fff2fff6ffff0000",
    56 => x"ffeefffcfffe0000",
    57 => x"fff1fffdfffe0000",
    58 => x"fff3fff3ffff0000",
    59 => x"fffcfffd00010000",
    60 => x"0005fff8ffff0000",
    61 => x"fffffffd00000000",
    62 => x"00050008ffff0000",
    63 => x"00170000ffff0000",
    64 => x"fff00000fffc0000",
    65 => x"fff3000dffff0000",
    66 => x"fff3000dffff0000",
    67 => x"fff0000000020000",
    68 => x"fff3000dffff0000",
    69 => x"00050008ffff0000",
    70 => x"0005000000010000",
    71 => x"ffff000300000000",
    72 => x"fff8000000020000",
    73 => x"fffc000300010000",
    74 => x"ffff000300000000",
    75 => x"fffc000300010000",
    76 => x"fffc000300010000",
    77 => x"fffc000000040000",
    78 => x"ffff000300000000",
    79 => x"0001000000040000",
    80 => x"00050008ffff0000",
    81 => x"000c0008ffff0000",
    82 => x"fff10003fffe0000",
    83 => x"fff1000300010000",
    84 => x"fff10003fffe0000",
    85 => x"fff2000affff0000",
    86 => x"fff2000affff0000",
    87 => x"fff1000300010000",
    88 => x"fff0000000020000",
    89 => x"fff1000300010000",
    90 => x"fff2000affff0000",
    91 => x"fff3000dffff0000",
    92 => x"fff10003fffe0000",
    93 => x"fff00000fffc0000",
    94 => x"ffee0004fffe0000",
    95 => x"ffee000400010000",
    96 => x"ffee0004fffe0000",
    97 => x"ffef000affff0000",
    98 => x"ffef000affff0000",
    99 => x"ffee000400010000",
    100 => x"fff1000300010000",
    101 => x"ffee000400010000",
    102 => x"ffef000affff0000",
    103 => x"fff2000affff0000",
    104 => x"ffee0004fffe0000",
    105 => x"fff10003fffe0000",
    106 => x"fff3000dffff0000",
    107 => x"fffc000300010000",
    108 => x"00050008ffff0000",
    109 => x"ffff000300000000",
    110 => x"ffffffffffffffff",
    111 => x"ffffffffffffffff",

    122 => x"fffaffee00160000",
    123 => x"fff8ffe900000000",
    124 => x"fff8ffe900000000",
    125 => x"0010fff6000c0000",
    126 => x"0010fff6000c0000",
    127 => x"fffaffee00160000",
    128 => x"0010fff6fff40000",
    129 => x"0010fff6000c0000",
    130 => x"fff8ffe900000000",
    131 => x"0010fff6fff40000",
    132 => x"ffeefffb00000000",
    133 => x"fff8ffe900000000",
    134 => x"fffaffee00160000",
    135 => x"ffeefffb00000000",
    136 => x"fffffff5ffec0000",
    137 => x"fff8ffe900000000",
    138 => x"ffeefffb00000000",
    139 => x"fffffff5ffec0000",
    140 => x"fffffff5ffec0000",
    141 => x"0010fff6fff40000",
    142 => x"0014000a00000000",
    143 => x"0010fff6000c0000",
    144 => x"0010fff6fff40000",
    145 => x"0014000a00000000",
    146 => x"0006000a00130000",
    147 => x"fffaffee00160000",
    148 => x"0010fff6000c0000",
    149 => x"0006000a00130000",
    150 => x"fff0000a000c0000",
    151 => x"ffeefffb00000000",
    152 => x"fffaffee00160000",
    153 => x"fff0000a000c0000",
    154 => x"ffec0007fff00000",
    155 => x"fffffff5ffec0000",
    156 => x"ffeefffb00000000",
    157 => x"ffec0007fff00000",
    158 => x"0006000affed0000",
    159 => x"0010fff6fff40000",
    160 => x"fffffff5ffec0000",
    161 => x"0006000affed0000",
    162 => x"0014000a00000000",
    163 => x"0006000a00130000",
    164 => x"0006000a00130000",
    165 => x"fff0000a000c0000",
    166 => x"fff0000a000c0000",
    167 => x"ffec0007fff00000",
    168 => x"ffec0007fff00000",
    169 => x"0006000affed0000",
    170 => x"0006000affed0000",
    171 => x"0014000a00000000",
    172 => x"0002001300060000",
    173 => x"0006000a00130000",
    174 => x"0014000a00000000",
    175 => x"0002001300060000",
    176 => x"0002001300060000",
    177 => x"fff0000a000c0000",
    178 => x"0002001300060000",
    179 => x"ffec0007fff00000",
    180 => x"0002001300060000",
    181 => x"0006000affed0000",
    182 => x"ffffffffffffffff",
    183 => x"ffffffffffffffff",



    --Start of asteroid
    190 => x"fffd0011ffef0000",
    191 => x"00020012ffed0000",
    192 => x"0003fff0fff40000",
    193 => x"0005fffefff20000",
    194 => x"ffff0010ffef0000",
    195 => x"00070010fff20000",
    196 => x"fffefffeffef0000",
    197 => x"fff8fffefff20000",
    198 => x"00070010fff20000",
    199 => x"000c0010fffe0000",
    200 => x"fff5fff0fffe0000",
    201 => x"fffefff0fffe0000",
    202 => x"fff80010fff20000",
    203 => x"ffff0010ffef0000",
    204 => x"0005fffefff20000",
    205 => x"fffefffeffef0000",
    206 => x"0006fff0fffe0000",
    207 => x"0004ffedfffe0000",
    208 => x"fff2fffefffe0000",
    209 => x"fff5fff0fffe0000",
    210 => x"fff8fffefff20000",
    211 => x"fff2fffefffe0000",
    212 => x"0006fff0fffe0000",
    213 => x"0003fff0fff40000",
    214 => x"fff5fff0fffe0000",
    215 => x"fff1ffecfffe0000",
    216 => x"fffefff0fffe0000",
    217 => x"0006fff0fffe0000",
    218 => x"fffeffedfff50000",
    219 => x"fff5fff0fffe0000",
    220 => x"fff8fffefff20000",
    221 => x"fffeffedfff50000",
    222 => x"000afffefffe0000",
    223 => x"0006fff0fffe0000",
    224 => x"0007001cfff50000",
    225 => x"00070010fff20000",
    226 => x"0004ffedfffe0000",
    227 => x"0003fff0fff40000",
    228 => x"fff1ffecfffe0000",
    229 => x"fffeffedfff50000",
    230 => x"00090028fff90000",
    231 => x"00090022fffe0000",
    232 => x"0002001cfff10000",
    233 => x"0007001cfff50000",
    234 => x"0007001cfff50000",
    235 => x"000b001cfffe0000",
    236 => x"fffc001cfff50000",
    237 => x"0002001cfff10000",
    238 => x"00030024fff60000",
    239 => x"00070024fff80000",
    240 => x"00070024fff80000",
    241 => x"00090022fffe0000",
    242 => x"00000025fff80000",
    243 => x"00030024fff60000",
    244 => x"0002001cfff10000",
    245 => x"00030024fff60000",
    246 => x"00070024fff80000",
    247 => x"0007001cfff50000",
    248 => x"fffc001cfff50000",
    249 => x"00000025fff80000",
    250 => x"00090022fffe0000",
    251 => x"000b001cfffe0000",
    252 => x"fff20010fffe0000",
    253 => x"fff2fffefffe0000",
    254 => x"fff7001cfffe0000",
    255 => x"fffd0025fffe0000",
    256 => x"00000025fff80000",
    257 => x"0006002afffa0000",
    258 => x"0006002afffa0000",
    259 => x"00070028fff80000",
    260 => x"fffd0025fffe0000",
    261 => x"0004002cfffe0000",
    262 => x"0009002afffa0000",
    263 => x"00090028fff90000",
    264 => x"0004002cfffe0000",
    265 => x"0009002bfffe0000",
    266 => x"0009002bfffe0000",
    267 => x"000d002afffe0000",
    268 => x"00070028fff80000",
    269 => x"00090028fff90000",
    270 => x"0006002afffa0000",
    271 => x"0009002afffa0000",
    272 => x"000d002afffe0000",
    273 => x"000d0028fffa0000",
    274 => x"000d002afffe0000",
    275 => x"0009002afffa0000",
    276 => x"00090028fff90000",
    277 => x"000d0028fffa0000",
    278 => x"00100028fffc0000",
    279 => x"00110027fffe0000",
    280 => x"000d0028fffa0000",
    281 => x"00100028fffc0000",
    282 => x"00070029fff90000",
    283 => x"00080029fff90000",
    284 => x"00080029fff90000",
    285 => x"00080029fff90000",
    286 => x"00080029fff90000",
    287 => x"00080029fff90000",
    288 => x"00070029fff90000",
    289 => x"00080029fff90000",
    290 => x"ffff0010ffef0000",
    291 => x"fffefffeffef0000",
    292 => x"00110027fffe0000",
    293 => x"00130028fffe0000",
    294 => x"00100029fffe0000",
    295 => x"00130028fffe0000",
    296 => x"00130028fffe0000",
    297 => x"00100028fffc0000",
    298 => x"fff80010fff20000",
    299 => x"fff8fffefff20000",
    300 => x"00100029fffe0000",
    301 => x"00100028fffc0000",
    302 => x"000d002afffe0000",
    303 => x"00100029fffe0000",
    304 => x"000d0028fffa0000",
    305 => x"000d0027fffe0000",
    306 => x"00070010fff20000",
    307 => x"0005fffefff20000",
    308 => x"00070028fff80000",
    309 => x"00030024fff60000",
    310 => x"fffd0011ffef0000",
    311 => x"fffffffdffeb0000",
    312 => x"fff20010fffe0000",
    313 => x"fff7001cfffe0000",
    314 => x"000afffefffe0000",
    315 => x"0005fffefff20000",
    316 => x"000c0010fffe0000",
    317 => x"000afffefffe0000",
    318 => x"000c0010fffe0000",
    319 => x"000b001cfffe0000",
    320 => x"fff20010fffe0000",
    321 => x"fff80010fff20000",
    322 => x"00020012ffed0000",
    323 => x"0002001cfff10000",
    324 => x"fffc001cfff50000",
    325 => x"fffd0011ffef0000",
    326 => x"fffffffdffeb0000",
    327 => x"0002fffcffe90000",
    328 => x"00060011ffef0000",
    329 => x"0007001cfff50000",
    330 => x"00020012ffed0000",
    331 => x"00060011ffef0000",
    332 => x"0002fffcffe90000",
    333 => x"00020012ffed0000",
    334 => x"00060011ffef0000",
    335 => x"0003fffeffeb0000",
    336 => x"fffc001cfff50000",
    337 => x"fff80010fff20000",
    338 => x"000d0027fffe0000",
    339 => x"00110027fffe0000",
    340 => x"0002fffcffe90000",
    341 => x"0003fffeffeb0000",
    342 => x"000d0027fffe0000",
    343 => x"00090022fffe0000",
    344 => x"00070028fff80000",
    345 => x"00070024fff80000",
    346 => x"ffff0010ffef0000",
    347 => x"0002001cfff10000",
    348 => x"fff7001cfffe0000",
    349 => x"fffc001cfff50000",
    350 => x"0004002cfffe0000",
    351 => x"0006002afffa0000",
    352 => x"fff1ffecfffe0000",
    353 => x"0004ffedfffe0000",
    354 => x"fffefff0fffe0000",
    355 => x"0004ffedfffe0000",
    356 => x"fffd0025fffe0000",
    357 => x"00000025fff80000",
    358 => x"0009002bfffe0000",
    359 => x"0009002afffa0000",
    360 => x"0004ffedfffe0000",
    361 => x"fffeffedfff50000",
    362 => x"0003fff0fff40000",
    363 => x"fffeffedfff50000",
    364 => x"fffefffeffef0000",
    365 => x"fffeffedfff50000",
    366 => x"fffd0011000c0000",
    367 => x"00020012000f0000",
    368 => x"0003fff000080000",
    369 => x"0005fffe000a0000",
    370 => x"ffff0010000d0000",
    371 => x"00070010000a0000",
    372 => x"fffefffe000d0000",
    373 => x"fff8fffe000a0000",
    374 => x"00070010000a0000",
    375 => x"000c0010fffe0000",
    376 => x"fff80010000a0000",
    377 => x"ffff0010000d0000",
    378 => x"0005fffe000a0000",
    379 => x"fffefffe000d0000",
    380 => x"fff8fffe000a0000",
    381 => x"fff2fffefffe0000",
    382 => x"0006fff0fffe0000",
    383 => x"0003fff000080000",
    384 => x"fffeffed00060000",
    385 => x"fff5fff0fffe0000",
    386 => x"fff8fffe000a0000",
    387 => x"fffeffed00060000",
    388 => x"0007001c00070000",
    389 => x"00070010000a0000",
    390 => x"0004ffedfffe0000",
    391 => x"0003fff000080000",
    392 => x"fff1ffecfffe0000",
    393 => x"fffeffed00060000",
    394 => x"0009002800030000",
    395 => x"00090022fffe0000",
    396 => x"0002001c000a0000",
    397 => x"0007001c00070000",
    398 => x"0007001c00070000",
    399 => x"000b001cfffe0000",
    400 => x"fffc001c00070000",
    401 => x"0002001c000a0000",
    402 => x"0003002400050000",
    403 => x"0007002400040000",
    404 => x"0007002400040000",
    405 => x"00090022fffe0000",
    406 => x"0000002500030000",
    407 => x"0003002400050000",
    408 => x"0002001c000a0000",
    409 => x"0003002400050000",
    410 => x"0007002400040000",
    411 => x"0007001c00070000",
    412 => x"fffc001c00070000",
    413 => x"0000002500030000",
    414 => x"0000002500030000",
    415 => x"0006002a00020000",
    416 => x"0006002a00020000",
    417 => x"0007002800040000",
    418 => x"0009002a00020000",
    419 => x"0009002800030000",
    420 => x"0007002800040000",
    421 => x"0009002800030000",
    422 => x"0006002a00020000",
    423 => x"0009002a00020000",
    424 => x"000d002afffe0000",
    425 => x"000d002800020000",
    426 => x"000d002afffe0000",
    427 => x"0009002a00020000",
    428 => x"0009002800030000",
    429 => x"000d002800020000",
    430 => x"0010002800000000",
    431 => x"00110027fffe0000",
    432 => x"000d002800020000",
    433 => x"0010002800000000",
    434 => x"0007002900030000",
    435 => x"0008002900030000",
    436 => x"0008002900030000",
    437 => x"0008002900030000",
    438 => x"0008002900030000",
    439 => x"0008002900030000",
    440 => x"0007002900030000",
    441 => x"0008002900030000",
    442 => x"ffff0010000d0000",
    443 => x"fffefffe000d0000",
    444 => x"00130028fffe0000",
    445 => x"0010002800000000",
    446 => x"fff80010000a0000",
    447 => x"fff8fffe000a0000",
    448 => x"00100029fffe0000",
    449 => x"0010002800000000",
    450 => x"000d002800020000",
    451 => x"000d0027fffe0000",
    452 => x"00070010000a0000",
    453 => x"0005fffe000a0000",
    454 => x"0007002800040000",
    455 => x"0003002400050000",
    456 => x"fffd0011000c0000",
    457 => x"fffffffd00110000",
    458 => x"000afffefffe0000",
    459 => x"0005fffe000a0000",
    460 => x"fff20010fffe0000",
    461 => x"fff80010000a0000",
    462 => x"00020012000f0000",
    463 => x"0002001c000a0000",
    464 => x"fffc001c00070000",
    465 => x"fffd0011000c0000",
    466 => x"fffffffd00110000",
    467 => x"0002fffc00120000",
    468 => x"00060011000d0000",
    469 => x"0007001c00070000",
    470 => x"00020012000f0000",
    471 => x"00060011000d0000",
    472 => x"0002fffc00120000",
    473 => x"00020012000f0000",
    474 => x"00060011000d0000",
    475 => x"0003fffe00110000",
    476 => x"fffc001c00070000",
    477 => x"fff80010000a0000",
    478 => x"0002fffc00120000",
    479 => x"0003fffe00110000",
    480 => x"0007002800040000",
    481 => x"0007002400040000",
    482 => x"ffff0010000d0000",
    483 => x"0002001c000a0000",
    484 => x"fff7001cfffe0000",
    485 => x"fffc001c00070000",
    486 => x"0004002cfffe0000",
    487 => x"0006002a00020000",
    488 => x"fffd0025fffe0000",
    489 => x"0000002500030000",
    490 => x"0009002bfffe0000",
    491 => x"0009002a00020000",
    492 => x"0004ffedfffe0000",
    493 => x"fffeffed00060000",
    494 => x"0003fff000080000",
    495 => x"fffeffed00060000",
    496 => x"fffefffe000d0000",
    497 => x"fffeffed00060000",
    498 => x"ffffffffffffffff",
    499 => x"ffffffffffffffff",



    508 => x"0000000000000000",
    509 => x"000f000000000000",
    510 => x"ffffffffffffffff",
    511 => x"ffffffffffffffff",
        others => (others => '0'));

begin

PROCESS(clk)
BEGIN
  if (rising_edge(clk)) then
    -- synkron skrivning/läsning port 1
    read_data <= ram(to_integer(read_addr));
  end if;
END PROCESS;

end Behavioral;
