
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Vector;

--Constants
package GPU_Info is
    --TODO: Optimse the size of obj addr and model addr
    --The length of the addresses and data in the object memory
    constant OBJ_ADDR_SIZE: positive := 12;
    constant OBJ_DATA_SIZE: positive := Vector.MEMORY_SIZE;

    subtype ObjAddr_t is unsigned(OBJ_ADDR_SIZE - 1 downto 0);
    subtype ObjData_t is std_logic_vector(OBJ_DATA_SIZE - 1 downto 0);

    constant MODEL_ADDR_SIZE: positive := 9;

    subtype ModelAddr_t is unsigned(MODEL_ADDR_SIZE - 1 downto 0);
    subtype ModelData_t is Vector.InMemory_t;
end package;

library IEEE;

use IEEE.Numeric_std.all;
use IEEE.std_logic_1164.all;

use work.Vector;
use work.GPU_Info;

entity ModelMem is
port (
        clk : in std_logic;
        -- port 1
        read_addr : in GPU_Info.ModelAddr_t;
        read_data : out GPU_Info.ModelData_t
    );
end entity;

architecture Behavioral of ModelMem is

-- Deklaration av ett dubbelportat block-RAM
-- med 2048 adresser av 8 bitars bredd.
type ram_t is array (0 to 4095) of Vector.InMemory_t;

    -- Nollställ alla bitar på alla adresser
    signal ram : ram_t := (
    0 => x"000e0000fffd0000",
    1 => x"000e000000020000",
    2 => x"ffeb000000000000",
    3 => x"000e0000fffd0000",
    4 => x"fffb000700000000",
    5 => x"ffeb000000000000",
    6 => x"fffc000000010000",
    7 => x"ffeb000000000000",
    8 => x"000e0000fffd0000",
    9 => x"000c000c00000000",
    10 => x"000c000c00000000",
    11 => x"000e000000020000",
    12 => x"000c000c00000000",
    13 => x"fffb000700000000",
    14 => x"000e000000020000",
    15 => x"0007000000020000",
    16 => x"0000000000030000",
    17 => x"fffc000000010000",
    18 => x"fffc000000010000",
    19 => x"0001000300000000",
    20 => x"0007000000020000",
    21 => x"0004000300010000",
    22 => x"0001000300000000",
    23 => x"0004000300010000",
    24 => x"0007000000020000",
    25 => x"0004000000040000",
    26 => x"0004000000040000",
    27 => x"0000000000030000",
    28 => x"0004000300010000",
    29 => x"0004000000040000",
    30 => x"0001000300000000",
    31 => x"0000000000030000",
    32 => x"fffb000700000000",
    33 => x"fff5000700000000",
    34 => x"000e0003fffe0000",
    35 => x"000e000300010000",
    36 => x"000e0003fffe0000",
    37 => x"000d000900000000",
    38 => x"000d000900000000",
    39 => x"000e000300010000",
    40 => x"000e000000020000",
    41 => x"000e000300010000",
    42 => x"000d000900000000",
    43 => x"000c000c00000000",
    44 => x"000e0003fffe0000",
    45 => x"000e0000fffd0000",
    46 => x"00100003fffe0000",
    47 => x"0010000300010000",
    48 => x"00100003fffe0000",
    49 => x"000f000900000000",
    50 => x"000f000900000000",
    51 => x"0010000300010000",
    52 => x"000e000300010000",
    53 => x"0010000300010000",
    54 => x"000f000900000000",
    55 => x"000d000900000000",
    56 => x"00100003fffe0000",
    57 => x"000e0003fffe0000",
    58 => x"000c000c00000000",
    59 => x"0004000300010000",
    60 => x"fffb000700000000",
    61 => x"0001000300000000",
    62 => x"fffbfff900000000",
    63 => x"ffeb000000000000",
    64 => x"000e0000fffd0000",
    65 => x"000cfff400000000",
    66 => x"000cfff400000000",
    67 => x"000e000000020000",
    68 => x"000cfff400000000",
    69 => x"fffbfff900000000",
    70 => x"fffc000000010000",
    71 => x"0001fffd00000000",
    72 => x"0007000000020000",
    73 => x"0004fffd00010000",
    74 => x"0001fffd00000000",
    75 => x"0004fffd00010000",
    76 => x"0004fffd00010000",
    77 => x"0004000000040000",
    78 => x"0001fffd00000000",
    79 => x"0000000000030000",
    80 => x"fffbfff900000000",
    81 => x"fff5fff900000000",
    82 => x"000efffdfffe0000",
    83 => x"000efffd00010000",
    84 => x"000efffdfffe0000",
    85 => x"000dfff700000000",
    86 => x"000dfff700000000",
    87 => x"000efffd00010000",
    88 => x"000e000000020000",
    89 => x"000efffd00010000",
    90 => x"000dfff700000000",
    91 => x"000cfff400000000",
    92 => x"000efffdfffe0000",
    93 => x"000e0000fffd0000",
    94 => x"0010fffdfffe0000",
    95 => x"0010fffd00010000",
    96 => x"0010fffdfffe0000",
    97 => x"000ffff700000000",
    98 => x"000ffff700000000",
    99 => x"0010fffd00010000",
    100 => x"000efffd00010000",
    101 => x"0010fffd00010000",
    102 => x"000ffff700000000",
    103 => x"000dfff700000000",
    104 => x"0010fffdfffe0000",
    105 => x"000efffdfffe0000",
    106 => x"000cfff400000000",
    107 => x"0004fffd00010000",
    108 => x"fffbfff900000000",
    109 => x"0001fffd00000000",
    110 => x"ffffffffffffffff",
    111 => x"ffffffffffffffff",

    --Start of asteroid
    122 => x"fffaffee00160000",
    123 => x"fff8ffe900000000",
    124 => x"fff8ffe900000000",
    125 => x"0010fff6000c0000",
    126 => x"0010fff6000c0000",
    127 => x"fffaffee00160000",
    128 => x"0010fff6fff40000",
    129 => x"0010fff6000c0000",
    130 => x"fff8ffe900000000",
    131 => x"0010fff6fff40000",
    132 => x"ffeefffb00000000",
    133 => x"fff8ffe900000000",
    134 => x"fffaffee00160000",
    135 => x"ffeefffb00000000",
    136 => x"fffffff5ffec0000",
    137 => x"fff8ffe900000000",
    138 => x"ffeefffb00000000",
    139 => x"fffffff5ffec0000",
    140 => x"fffffff5ffec0000",
    141 => x"0010fff6fff40000",
    142 => x"0014000a00000000",
    143 => x"0010fff6000c0000",
    144 => x"0010fff6fff40000",
    145 => x"0014000a00000000",
    146 => x"0006000a00130000",
    147 => x"fffaffee00160000",
    148 => x"0010fff6000c0000",
    149 => x"0006000a00130000",
    150 => x"fff0000a000c0000",
    151 => x"ffeefffb00000000",
    152 => x"fffaffee00160000",
    153 => x"fff0000a000c0000",
    154 => x"ffec0007fff00000",
    155 => x"fffffff5ffec0000",
    156 => x"ffeefffb00000000",
    157 => x"ffec0007fff00000",
    158 => x"0006000affed0000",
    159 => x"0010fff6fff40000",
    160 => x"fffffff5ffec0000",
    161 => x"0006000affed0000",
    162 => x"0014000a00000000",
    163 => x"0006000a00130000",
    164 => x"0006000a00130000",
    165 => x"fff0000a000c0000",
    166 => x"fff0000a000c0000",
    167 => x"ffec0007fff00000",
    168 => x"ffec0007fff00000",
    169 => x"0006000affed0000",
    170 => x"0006000affed0000",
    171 => x"0014000a00000000",
    172 => x"0002001300060000",
    173 => x"0006000a00130000",
    174 => x"0014000a00000000",
    175 => x"0002001300060000",
    176 => x"0002001300060000",
    177 => x"fff0000a000c0000",
    178 => x"0002001300060000",
    179 => x"ffec0007fff00000",
    180 => x"0002001300060000",
    181 => x"0006000affed0000",
    182 => x"ffffffffffffffff",
    183 => x"ffffffffffffffff",

    190 => x"0040001400280000",
    191 => x"0035001400310000",
    192 => x"0035001400310000",
    193 => x"0032000b00320000",
    194 => x"0032000b00320000",
    195 => x"0039000300290000",
    196 => x"0039000300290000",
    197 => x"0040001400280000",
    198 => x"ffc0001400280000",
    199 => x"ffc7000300290000",
    200 => x"ffc7000300290000",
    201 => x"ffce000b00320000",
    202 => x"ffce000b00320000",
    203 => x"ffcb001400310000",
    204 => x"ffcb001400310000",
    205 => x"ffc0001400280000",
    206 => x"00470014001b0000",
    207 => x"0040001400280000",
    208 => x"0039000300290000",
    209 => x"003effff001d0000",
    210 => x"003effff001d0000",
    211 => x"00470014001b0000",
    212 => x"ffb90014001b0000",
    213 => x"ffc2ffff001d0000",
    214 => x"ffc2ffff001d0000",
    215 => x"ffc7000300290000",
    216 => x"ffc0001400280000",
    217 => x"ffb90014001b0000",
    218 => x"0039000300290000",
    219 => x"0028fffc002d0000",
    220 => x"0028fffc002d0000",
    221 => x"0028fff600210000",
    222 => x"0028fff600210000",
    223 => x"003effff001d0000",
    224 => x"ffc2ffff001d0000",
    225 => x"ffd8fff600210000",
    226 => x"ffd8fff600210000",
    227 => x"ffd8fffc002d0000",
    228 => x"ffd8fffc002d0000",
    229 => x"ffc7000300290000",
    230 => x"0032000b00320000",
    231 => x"0028000700340000",
    232 => x"0028000700340000",
    233 => x"0028fffc002d0000",
    234 => x"ffd8fffc002d0000",
    235 => x"ffd8000700340000",
    236 => x"ffd8000700340000",
    237 => x"ffce000b00320000",
    238 => x"0028000700340000",
    239 => x"001f000b00360000",
    240 => x"001f000b00360000",
    241 => x"0017000300300000",
    242 => x"0017000300300000",
    243 => x"0028fffc002d0000",
    244 => x"ffd8fffc002d0000",
    245 => x"ffe9000300300000",
    246 => x"ffe9000300300000",
    247 => x"ffe1000b00360000",
    248 => x"ffe1000b00360000",
    249 => x"ffd8000700340000",
    250 => x"0017000300300000",
    251 => x"0012ffff00250000",
    252 => x"0012ffff00250000",
    253 => x"0028fff600210000",
    254 => x"ffd8fff600210000",
    255 => x"ffeeffff00250000",
    256 => x"ffeeffff00250000",
    257 => x"ffe9000300300000",
    258 => x"0017000300300000",
    259 => x"0010001400300000",
    260 => x"0010001400300000",
    261 => x"0009001400260000",
    262 => x"0009001400260000",
    263 => x"0012ffff00250000",
    264 => x"ffeeffff00250000",
    265 => x"fff7001400260000",
    266 => x"fff7001400260000",
    267 => x"fff0001400300000",
    268 => x"fff0001400300000",
    269 => x"ffe9000300300000",
    270 => x"001f000b00360000",
    271 => x"001c001400360000",
    272 => x"001c001400360000",
    273 => x"0010001400300000",
    274 => x"fff0001400300000",
    275 => x"ffe4001400360000",
    276 => x"ffe4001400360000",
    277 => x"ffe1000b00360000",
    278 => x"001c001400360000",
    279 => x"001f001e00360000",
    280 => x"001f001e00360000",
    281 => x"0017002500300000",
    282 => x"0017002500300000",
    283 => x"0010001400300000",
    284 => x"fff0001400300000",
    285 => x"ffe9002500300000",
    286 => x"ffe9002500300000",
    287 => x"ffe1001e00360000",
    288 => x"ffe1001e00360000",
    289 => x"ffe4001400360000",
    290 => x"0017002500300000",
    291 => x"0012002a00250000",
    292 => x"0012002a00250000",
    293 => x"0009001400260000",
    294 => x"fff7001400260000",
    295 => x"ffee002a00250000",
    296 => x"ffee002a00250000",
    297 => x"ffe9002500300000",
    298 => x"0017002500300000",
    299 => x"0028002c002d0000",
    300 => x"0028002c002d0000",
    301 => x"0028003300210000",
    302 => x"0028003300210000",
    303 => x"0012002a00250000",
    304 => x"ffee002a00250000",
    305 => x"ffd8003300210000",
    306 => x"ffd8003300210000",
    307 => x"ffd8002c002d0000",
    308 => x"ffd8002c002d0000",
    309 => x"ffe9002500300000",
    310 => x"001f001e00360000",
    311 => x"0028002100340000",
    312 => x"0028002100340000",
    313 => x"0028002c002d0000",
    314 => x"ffd8002c002d0000",
    315 => x"ffd8002100340000",
    316 => x"ffd8002100340000",
    317 => x"ffe1001e00360000",
    318 => x"0028002100340000",
    319 => x"0032001e00320000",
    320 => x"0032001e00320000",
    321 => x"0039002500290000",
    322 => x"0039002500290000",
    323 => x"0028002c002d0000",
    324 => x"ffd8002c002d0000",
    325 => x"ffc7002500290000",
    326 => x"ffc7002500290000",
    327 => x"ffce001e00320000",
    328 => x"ffce001e00320000",
    329 => x"ffd8002100340000",
    330 => x"0039002500290000",
    331 => x"003e002a001d0000",
    332 => x"003e002a001d0000",
    333 => x"0028003300210000",
    334 => x"ffd8003300210000",
    335 => x"ffc2002a001d0000",
    336 => x"ffc2002a001d0000",
    337 => x"ffc7002500290000",
    338 => x"0039002500290000",
    339 => x"0040001400280000",
    340 => x"00470014001b0000",
    341 => x"003e002a001d0000",
    342 => x"ffc2002a001d0000",
    343 => x"ffb90014001b0000",
    344 => x"ffc0001400280000",
    345 => x"ffc7002500290000",
    346 => x"0032001e00320000",
    347 => x"0035001400310000",
    348 => x"ffcb001400310000",
    349 => x"ffce001e00320000",
    350 => x"0036001400330000",
    351 => x"0035001400310000",
    352 => x"0032001e00320000",
    353 => x"0033001f00340000",
    354 => x"0033001f00340000",
    355 => x"0036001400330000",
    356 => x"ffca001400330000",
    357 => x"ffcd001f00340000",
    358 => x"ffcd001f00340000",
    359 => x"ffce001e00320000",
    360 => x"ffcb001400310000",
    361 => x"ffca001400330000",
    362 => x"0028002100340000",
    363 => x"0028002300370000",
    364 => x"0028002300370000",
    365 => x"0033001f00340000",
    366 => x"ffcd001f00340000",
    367 => x"ffd8002300370000",
    368 => x"ffd8002300370000",
    369 => x"ffd8002100340000",
    370 => x"001f001e00360000",
    371 => x"001e001f00380000",
    372 => x"001e001f00380000",
    373 => x"0028002300370000",
    374 => x"ffd8002300370000",
    375 => x"ffe2001f00380000",
    376 => x"ffe2001f00380000",
    377 => x"ffe1001e00360000",
    378 => x"001c001400360000",
    379 => x"001a001400380000",
    380 => x"001a001400380000",
    381 => x"001e001f00380000",
    382 => x"ffe2001f00380000",
    383 => x"ffe6001400380000",
    384 => x"ffe6001400380000",
    385 => x"ffe4001400360000",
    386 => x"001f000b00360000",
    387 => x"001e000a00380000",
    388 => x"001e000a00380000",
    389 => x"001a001400380000",
    390 => x"ffe6001400380000",
    391 => x"ffe2000a00380000",
    392 => x"ffe2000a00380000",
    393 => x"ffe1000b00360000",
    394 => x"0028000700340000",
    395 => x"0028000600370000",
    396 => x"0028000600370000",
    397 => x"001e000a00380000",
    398 => x"ffe2000a00380000",
    399 => x"ffd8000600370000",
    400 => x"ffd8000600370000",
    401 => x"ffd8000700340000",
    402 => x"0032000b00320000",
    403 => x"0033000a00340000",
    404 => x"0033000a00340000",
    405 => x"0028000600370000",
    406 => x"ffd8000600370000",
    407 => x"ffcd000a00340000",
    408 => x"ffcd000a00340000",
    409 => x"ffce000b00320000",
    410 => x"0036001400330000",
    411 => x"0033000a00340000",
    412 => x"ffcd000a00340000",
    413 => x"ffca001400330000",
    414 => x"0036001400330000",
    415 => x"0028001400390000",
    416 => x"0028001400390000",
    417 => x"0033000a00340000",
    418 => x"ffd8001400390000",
    419 => x"ffca001400330000",
    420 => x"ffcd000a00340000",
    421 => x"ffd8001400390000",
    422 => x"0028001400390000",
    423 => x"0028000600370000",
    424 => x"ffd8000600370000",
    425 => x"ffd8001400390000",
    426 => x"0028001400390000",
    427 => x"001e000a00380000",
    428 => x"ffe2000a00380000",
    429 => x"ffd8001400390000",
    430 => x"0028001400390000",
    431 => x"001a001400380000",
    432 => x"ffe6001400380000",
    433 => x"ffd8001400390000",
    434 => x"0028001400390000",
    435 => x"001e001f00380000",
    436 => x"ffe2001f00380000",
    437 => x"ffd8001400390000",
    438 => x"0028001400390000",
    439 => x"0028002300370000",
    440 => x"ffd8002300370000",
    441 => x"ffd8001400390000",
    442 => x"0028001400390000",
    443 => x"0033001f00340000",
    444 => x"ffcd001f00340000",
    445 => x"ffd8001400390000",
    446 => x"0000ff88001d0000",
    447 => x"0014ff8a001a0000",
    448 => x"0014ff8a001a0000",
    449 => x"0013ff8f00230000",
    450 => x"0013ff8f00230000",
    451 => x"0000ff8d00240000",
    452 => x"0000ff8d00240000",
    453 => x"0000ff88001d0000",
    454 => x"0000ff8d00240000",
    455 => x"ffedff8f00230000",
    456 => x"ffedff8f00230000",
    457 => x"ffecff8a001a0000",
    458 => x"ffecff8a001a0000",
    459 => x"0000ff88001d0000",
    460 => x"0014ff8a001a0000",
    461 => x"0025ff8d00170000",
    462 => x"0025ff8d00170000",
    463 => x"001bff9000230000",
    464 => x"001bff9000230000",
    465 => x"0013ff8f00230000",
    466 => x"ffedff8f00230000",
    467 => x"ffe5ff9000230000",
    468 => x"ffe5ff9000230000",
    469 => x"ffdbff8d00170000",
    470 => x"ffdbff8d00170000",
    471 => x"ffecff8a001a0000",
    472 => x"0025ff8d00170000",
    473 => x"002aff9300180000",
    474 => x"002aff9300180000",
    475 => x"001eff9b00270000",
    476 => x"001eff9b00270000",
    477 => x"001bff9000230000",
    478 => x"ffe5ff9000230000",
    479 => x"ffe2ff9b00270000",
    480 => x"ffe2ff9b00270000",
    481 => x"ffd6ff9300180000",
    482 => x"ffd6ff9300180000",
    483 => x"ffdbff8d00170000",
    484 => x"002aff9300180000",
    485 => x"0028ffa9001c0000",
    486 => x"0028ffa9001c0000",
    487 => x"001cffa800290000",
    488 => x"001cffa800290000",
    489 => x"001eff9b00270000",
    490 => x"ffe2ff9b00270000",
    491 => x"ffe4ffa800290000",
    492 => x"ffe4ffa800290000",
    493 => x"ffd8ffa9001c0000",
    494 => x"ffd8ffa9001c0000",
    495 => x"ffd6ff9300180000",
    496 => x"0028ffa9001c0000",
    497 => x"0024ffc7001c0000",
    498 => x"0024ffc7001c0000",
    499 => x"0018ffc6002c0000",
    500 => x"0018ffc6002c0000",
    501 => x"001cffa800290000",
    502 => x"ffe4ffa800290000",
    503 => x"ffe8ffc6002c0000",
    504 => x"ffe8ffc6002c0000",
    505 => x"ffdcffc7001c0000",
    506 => x"ffdcffc7001c0000",
    507 => x"ffd8ffa9001c0000",
    508 => x"000effed00380000",
    509 => x"0017ffe3001b0000",
    510 => x"0017ffe3001b0000",
    511 => x"0032ffe800180000",
    512 => x"0032ffe800180000",
    513 => x"002dfff300280000",
    514 => x"002dfff300280000",
    515 => x"000effed00380000",
    516 => x"fff2ffed00380000",
    517 => x"ffd3fff300280000",
    518 => x"ffd3fff300280000",
    519 => x"ffceffe800180000",
    520 => x"ffceffe800180000",
    521 => x"ffe9ffe3001b0000",
    522 => x"ffe9ffe3001b0000",
    523 => x"fff2ffed00380000",
    524 => x"0032ffe800180000",
    525 => x"0048fff400180000",
    526 => x"0048fff400180000",
    527 => x"0046ffff00220000",
    528 => x"0046ffff00220000",
    529 => x"002dfff300280000",
    530 => x"ffd3fff300280000",
    531 => x"ffbaffff00220000",
    532 => x"ffbaffff00220000",
    533 => x"ffb8fff400180000",
    534 => x"ffb8fff400180000",
    535 => x"ffceffe800180000",
    536 => x"0048fff400180000",
    537 => x"005e0009000e0000",
    538 => x"005e0009000e0000",
    539 => x"0053000f00200000",
    540 => x"0053000f00200000",
    541 => x"0046ffff00220000",
    542 => x"ffbaffff00220000",
    543 => x"ffad000f00200000",
    544 => x"ffad000f00200000",
    545 => x"ffa20009000e0000",
    546 => x"ffa20009000e0000",
    547 => x"ffb8fff400180000",
    548 => x"005e0009000e0000",
    549 => x"00620029001f0000",
    550 => x"00620029001f0000",
    551 => x"0054002300260000",
    552 => x"0054002300260000",
    553 => x"0053000f00200000",
    554 => x"ffad000f00200000",
    555 => x"ffac002300260000",
    556 => x"ffac002300260000",
    557 => x"ff9e0029001f0000",
    558 => x"ff9e0029001f0000",
    559 => x"ffa20009000e0000",
    560 => x"00620029001f0000",
    561 => x"0051002f00220000",
    562 => x"0051002f00220000",
    563 => x"004e0027002e0000",
    564 => x"004e0027002e0000",
    565 => x"0054002300260000",
    566 => x"ffac002300260000",
    567 => x"ffb20027002e0000",
    568 => x"ffb20027002e0000",
    569 => x"ffaf002f00220000",
    570 => x"ffaf002f00220000",
    571 => x"ff9e0029001f0000",
    572 => x"0051002f00220000",
    573 => x"0038003d00290000",
    574 => x"0038003d00290000",
    575 => x"0032003700360000",
    576 => x"0032003700360000",
    577 => x"004e0027002e0000",
    578 => x"ffb20027002e0000",
    579 => x"ffce003700360000",
    580 => x"ffce003700360000",
    581 => x"ffc8003d00290000",
    582 => x"ffc8003d00290000",
    583 => x"ffaf002f00220000",
    584 => x"0038003d00290000",
    585 => x"0024004e002f0000",
    586 => x"0024004e002f0000",
    587 => x"00240041003a0000",
    588 => x"00240041003a0000",
    589 => x"0032003700360000",
    590 => x"ffce003700360000",
    591 => x"ffdc0041003a0000",
    592 => x"ffdc0041003a0000",
    593 => x"ffdc004e002f0000",
    594 => x"ffdc004e002f0000",
    595 => x"ffc8003d00290000",
    596 => x"0024004e002f0000",
    597 => x"0012004a00310000",
    598 => x"0012004a00310000",
    599 => x"0017003f003c0000",
    600 => x"0017003f003c0000",
    601 => x"00240041003a0000",
    602 => x"ffdc0041003a0000",
    603 => x"ffe9003f003c0000",
    604 => x"ffe9003f003c0000",
    605 => x"ffee004a00310000",
    606 => x"ffee004a00310000",
    607 => x"ffdc004e002f0000",
    608 => x"0012004a00310000",
    609 => x"0007003000300000",
    610 => x"0007003000300000",
    611 => x"000c0029003b0000",
    612 => x"000c0029003b0000",
    613 => x"0017003f003c0000",
    614 => x"ffe9003f003c0000",
    615 => x"fff40029003b0000",
    616 => x"fff40029003b0000",
    617 => x"fff9003000300000",
    618 => x"fff9003000300000",
    619 => x"ffee004a00310000",
    620 => x"0007003000300000",
    621 => x"0000002900300000",
    622 => x"0000002900300000",
    623 => x"0000002000380000",
    624 => x"0000002000380000",
    625 => x"000c0029003b0000",
    626 => x"fff40029003b0000",
    627 => x"0000002000380000",
    628 => x"0000002900300000",
    629 => x"fff9003000300000",
    630 => x"000c0029003b0000",
    631 => x"0013002700330000",
    632 => x"0013002700330000",
    633 => x"001c002e00310000",
    634 => x"001c002e00310000",
    635 => x"0017003f003c0000",
    636 => x"ffe9003f003c0000",
    637 => x"ffe4002e00310000",
    638 => x"ffe4002e00310000",
    639 => x"ffed002700330000",
    640 => x"ffed002700330000",
    641 => x"fff40029003b0000",
    642 => x"001c002e00310000",
    643 => x"0025002f00300000",
    644 => x"0025002f00300000",
    645 => x"00240041003a0000",
    646 => x"ffdc0041003a0000",
    647 => x"ffdb002f00300000",
    648 => x"ffdb002f00300000",
    649 => x"ffe4002e00310000",
    650 => x"0025002f00300000",
    651 => x"0031002a002d0000",
    652 => x"0031002a002d0000",
    653 => x"0032003700360000",
    654 => x"ffce003700360000",
    655 => x"ffcf002a002d0000",
    656 => x"ffcf002a002d0000",
    657 => x"ffdb002f00300000",
    658 => x"0031002a002d0000",
    659 => x"0044002300270000",
    660 => x"0044002300270000",
    661 => x"004e0027002e0000",
    662 => x"ffb20027002e0000",
    663 => x"ffbc002300270000",
    664 => x"ffbc002300270000",
    665 => x"ffcf002a002d0000",
    666 => x"0044002300270000",
    667 => x"0049001a00250000",
    668 => x"0049001a00250000",
    669 => x"0054002300260000",
    670 => x"ffac002300260000",
    671 => x"ffb7001a00250000",
    672 => x"ffb7001a00250000",
    673 => x"ffbc002300270000",
    674 => x"0049001a00250000",
    675 => x"0047000e00250000",
    676 => x"0047000e00250000",
    677 => x"0053000f00200000",
    678 => x"ffad000f00200000",
    679 => x"ffb9000e00250000",
    680 => x"ffb9000e00250000",
    681 => x"ffb7001a00250000",
    682 => x"0047000e00250000",
    683 => x"0038ffff00280000",
    684 => x"0038ffff00280000",
    685 => x"0046ffff00220000",
    686 => x"ffbaffff00220000",
    687 => x"ffc8ffff00280000",
    688 => x"ffc8ffff00280000",
    689 => x"ffb9000e00250000",
    690 => x"0038ffff00280000",
    691 => x"002bfffa002b0000",
    692 => x"002bfffa002b0000",
    693 => x"002dfff300280000",
    694 => x"ffd3fff300280000",
    695 => x"ffd5fffa002b0000",
    696 => x"ffd5fffa002b0000",
    697 => x"ffc8ffff00280000",
    698 => x"002bfffa002b0000",
    699 => x"0017000300300000",
    700 => x"0017000300300000",
    701 => x"000effed00380000",
    702 => x"fff2ffed00380000",
    703 => x"ffe9000300300000",
    704 => x"ffe9000300300000",
    705 => x"ffd5fffa002b0000",
    706 => x"0017000300300000",
    707 => x"0013000800300000",
    708 => x"0013000800300000",
    709 => x"0000fffe002e0000",
    710 => x"0000fffe002e0000",
    711 => x"000effed00380000",
    712 => x"fff2ffed00380000",
    713 => x"0000fffe002e0000",
    714 => x"0000fffe002e0000",
    715 => x"ffed000800300000",
    716 => x"ffed000800300000",
    717 => x"ffe9000300300000",
    718 => x"000e001b00320000",
    719 => x"0013002700330000",
    720 => x"0000002000380000",
    721 => x"000e001b00320000",
    722 => x"fff2001b00320000",
    723 => x"0000002000380000",
    724 => x"ffed002700330000",
    725 => x"fff2001b00320000",
    726 => x"000f001000310000",
    727 => x"000e001b00320000",
    728 => x"0000002000380000",
    729 => x"0000001000320000",
    730 => x"0000001000320000",
    731 => x"000f001000310000",
    732 => x"fff1001000310000",
    733 => x"0000001000320000",
    734 => x"fff2001b00320000",
    735 => x"fff1001000310000",
    736 => x"0000001000320000",
    737 => x"0000fffe002e0000",
    738 => x"0013000800300000",
    739 => x"000f001000310000",
    740 => x"fff1001000310000",
    741 => x"ffed000800300000",
    742 => x"0013ff8f00230000",
    743 => x"0007ff94002a0000",
    744 => x"0007ff94002a0000",
    745 => x"0000ff9300290000",
    746 => x"0000ff9300290000",
    747 => x"0000ff8d00240000",
    748 => x"0000ff9300290000",
    749 => x"fff9ff94002a0000",
    750 => x"fff9ff94002a0000",
    751 => x"ffedff8f00230000",
    752 => x"001bff9000230000",
    753 => x"000dff99002c0000",
    754 => x"000dff99002c0000",
    755 => x"0007ff94002a0000",
    756 => x"fff9ff94002a0000",
    757 => x"fff3ff99002c0000",
    758 => x"fff3ff99002c0000",
    759 => x"ffe5ff9000230000",
    760 => x"001eff9b00270000",
    761 => x"000cffa7002f0000",
    762 => x"000cffa7002f0000",
    763 => x"000dff99002c0000",
    764 => x"fff3ff99002c0000",
    765 => x"fff4ffa7002f0000",
    766 => x"fff4ffa7002f0000",
    767 => x"ffe2ff9b00270000",
    768 => x"0018ffc6002c0000",
    769 => x"0009ffc600300000",
    770 => x"0009ffc600300000",
    771 => x"000dffaa002f0000",
    772 => x"000dffaa002f0000",
    773 => x"001cffa800290000",
    774 => x"ffe4ffa800290000",
    775 => x"fff3ffaa002f0000",
    776 => x"fff3ffaa002f0000",
    777 => x"fff7ffc600300000",
    778 => x"fff7ffc600300000",
    779 => x"ffe8ffc6002c0000",
    780 => x"000dffaa002f0000",
    781 => x"000cffa7002f0000",
    782 => x"fff4ffa7002f0000",
    783 => x"fff3ffaa002f0000",
    784 => x"0009ffc600300000",
    785 => x"000affd700300000",
    786 => x"000affd700300000",
    787 => x"0000ffd300300000",
    788 => x"0000ffd300300000",
    789 => x"0000ffc600300000",
    790 => x"0000ffc600300000",
    791 => x"0009ffc600300000",
    792 => x"fff7ffc600300000",
    793 => x"0000ffc600300000",
    794 => x"0000ffd300300000",
    795 => x"fff6ffd700300000",
    796 => x"fff6ffd700300000",
    797 => x"fff7ffc600300000",
    798 => x"0000ffab002f0000",
    799 => x"000dffaa002f0000",
    800 => x"0000ffc600300000",
    801 => x"0000ffab002f0000",
    802 => x"fff3ffaa002f0000",
    803 => x"0000ffab002f0000",
    804 => x"0000ffab002f0000",
    805 => x"0000ffa1002f0000",
    806 => x"0000ffa1002f0000",
    807 => x"000cffa7002f0000",
    808 => x"fff4ffa7002f0000",
    809 => x"0000ffa1002f0000",
    810 => x"000affd700300000",
    811 => x"000effdf00300000",
    812 => x"000effdf00300000",
    813 => x"000fffdf00360000",
    814 => x"000fffdf00360000",
    815 => x"000bffd900340000",
    816 => x"000bffd900340000",
    817 => x"000affd700300000",
    818 => x"fff6ffd700300000",
    819 => x"fff5ffd900340000",
    820 => x"fff5ffd900340000",
    821 => x"fff1ffdf00360000",
    822 => x"fff1ffdf00360000",
    823 => x"fff2ffdf00300000",
    824 => x"fff2ffdf00300000",
    825 => x"fff6ffd700300000",
    826 => x"000effdf00300000",
    827 => x"000cffe700300000",
    828 => x"000cffe700300000",
    829 => x"000cffe900340000",
    830 => x"000cffe900340000",
    831 => x"000fffdf00360000",
    832 => x"fff1ffdf00360000",
    833 => x"fff4ffe900340000",
    834 => x"fff4ffe900340000",
    835 => x"fff4ffe700300000",
    836 => x"fff4ffe700300000",
    837 => x"fff2ffdf00300000",
    838 => x"000cffe700300000",
    839 => x"0000ffe800300000",
    840 => x"0000ffe800300000",
    841 => x"0004ffea00340000",
    842 => x"0004ffea00340000",
    843 => x"000cffe900340000",
    844 => x"fff4ffe900340000",
    845 => x"fffcffea00340000",
    846 => x"fffcffea00340000",
    847 => x"0000ffe800300000",
    848 => x"0000ffe800300000",
    849 => x"fff4ffe700300000",
    850 => x"0000ffe800300000",
    851 => x"0000ffe200300000",
    852 => x"0000ffe200300000",
    853 => x"0000ffe300360000",
    854 => x"0000ffe300360000",
    855 => x"0004ffea00340000",
    856 => x"fffcffea00340000",
    857 => x"0000ffe300360000",
    858 => x"0000ffd400340000",
    859 => x"0000ffd300300000",
    860 => x"000bffd900340000",
    861 => x"0000ffd400340000",
    862 => x"0000ffd400340000",
    863 => x"fff5ffd900340000",
    864 => x"0000ffd700370000",
    865 => x"0000ffd400340000",
    866 => x"000bffd900340000",
    867 => x"0009ffdc00370000",
    868 => x"0009ffdc00370000",
    869 => x"0000ffd700370000",
    870 => x"0000ffd700370000",
    871 => x"fff7ffdc00370000",
    872 => x"fff7ffdc00370000",
    873 => x"fff5ffd900340000",
    874 => x"0000ffe300360000",
    875 => x"0000ffe100390000",
    876 => x"0000ffe100390000",
    877 => x"0005ffe700380000",
    878 => x"0005ffe700380000",
    879 => x"0004ffea00340000",
    880 => x"fffcffea00340000",
    881 => x"fffbffe700380000",
    882 => x"fffbffe700380000",
    883 => x"0000ffe100390000",
    884 => x"0005ffe700380000",
    885 => x"000bffe700380000",
    886 => x"000bffe700380000",
    887 => x"000cffe900340000",
    888 => x"fff4ffe900340000",
    889 => x"fff5ffe700380000",
    890 => x"fff5ffe700380000",
    891 => x"fffbffe700380000",
    892 => x"000bffe700380000",
    893 => x"000cffdf00390000",
    894 => x"000cffdf00390000",
    895 => x"000fffdf00360000",
    896 => x"fff1ffdf00360000",
    897 => x"fff4ffdf00390000",
    898 => x"fff4ffdf00390000",
    899 => x"fff5ffe700380000",
    900 => x"000cffdf00390000",
    901 => x"0009ffdc00370000",
    902 => x"fff7ffdc00370000",
    903 => x"fff4ffdf00390000",
    904 => x"0000ffe100390000",
    905 => x"000cffdf00390000",
    906 => x"fff4ffdf00390000",
    907 => x"0000ffe100390000",
    908 => x"0000ffe100390000",
    909 => x"0000ffd700370000",
    910 => x"0000fffe002e0000",
    911 => x"0000ffe800300000",
    912 => x"000cffe700300000",
    913 => x"000effed00380000",
    914 => x"fff2ffed00380000",
    915 => x"fff4ffe700300000",
    916 => x"000effdf00300000",
    917 => x"0013ffdd002c0000",
    918 => x"0013ffdd002c0000",
    919 => x"000effed00380000",
    920 => x"fff2ffed00380000",
    921 => x"ffedffdd002c0000",
    922 => x"ffedffdd002c0000",
    923 => x"fff2ffdf00300000",
    924 => x"000affd700300000",
    925 => x"0014ffd5002c0000",
    926 => x"0014ffd5002c0000",
    927 => x"0013ffdd002c0000",
    928 => x"ffedffdd002c0000",
    929 => x"ffecffd5002c0000",
    930 => x"ffecffd5002c0000",
    931 => x"fff6ffd700300000",
    932 => x"0018ffc6002c0000",
    933 => x"0014ffd5002c0000",
    934 => x"ffecffd5002c0000",
    935 => x"ffe8ffc6002c0000",
    936 => x"0024ffc7001c0000",
    937 => x"001dffd5001a0000",
    938 => x"001dffd5001a0000",
    939 => x"0014ffd5002c0000",
    940 => x"ffecffd5002c0000",
    941 => x"ffe3ffd5001a0000",
    942 => x"ffe3ffd5001a0000",
    943 => x"ffdcffc7001c0000",
    944 => x"001dffd5001a0000",
    945 => x"001bffdc001a0000",
    946 => x"001bffdc001a0000",
    947 => x"0013ffdd002c0000",
    948 => x"ffedffdd002c0000",
    949 => x"ffe5ffdc001a0000",
    950 => x"ffe5ffdc001a0000",
    951 => x"ffe3ffd5001a0000",
    952 => x"001bffdc001a0000",
    953 => x"0017ffe3001b0000",
    954 => x"ffe9ffe3001b0000",
    955 => x"ffe5ffdc001a0000",
    956 => x"000bffa4002e0000",
    957 => x"000cffa7002f0000",
    958 => x"0000ffa1002f0000",
    959 => x"0000ffa0002d0000",
    960 => x"0000ffa0002d0000",
    961 => x"000bffa4002e0000",
    962 => x"fff5ffa4002e0000",
    963 => x"0000ffa0002d0000",
    964 => x"fff4ffa7002f0000",
    965 => x"fff5ffa4002e0000",
    966 => x"000bff9b002c0000",
    967 => x"000dff99002c0000",
    968 => x"000bffa4002e0000",
    969 => x"000bff9b002c0000",
    970 => x"fff5ff9b002c0000",
    971 => x"fff5ffa4002e0000",
    972 => x"fff3ff99002c0000",
    973 => x"fff5ff9b002c0000",
    974 => x"0005ff9600290000",
    975 => x"0007ff94002a0000",
    976 => x"000bff9b002c0000",
    977 => x"0005ff9600290000",
    978 => x"fffbff9600290000",
    979 => x"fff5ff9b002c0000",
    980 => x"fff9ff94002a0000",
    981 => x"fffbff9600290000",
    982 => x"0000ff9500290000",
    983 => x"0000ff9300290000",
    984 => x"0005ff9600290000",
    985 => x"0000ff9500290000",
    986 => x"0000ff9500290000",
    987 => x"fffbff9600290000",
    988 => x"0000ff9700230000",
    989 => x"0000ff9500290000",
    990 => x"0005ff9600290000",
    991 => x"0005ff9700230000",
    992 => x"0005ff9700230000",
    993 => x"0000ff9700230000",
    994 => x"0000ff9700230000",
    995 => x"fffbff9700230000",
    996 => x"fffbff9700230000",
    997 => x"fffbff9600290000",
    998 => x"000bff9b002c0000",
    999 => x"000bff9c00240000",
    1000 => x"000bff9c00240000",
    1001 => x"0005ff9700230000",
    1002 => x"fffbff9700230000",
    1003 => x"fff5ff9c00240000",
    1004 => x"fff5ff9c00240000",
    1005 => x"fff5ff9b002c0000",
    1006 => x"000bffa4002e0000",
    1007 => x"000bffa300270000",
    1008 => x"000bffa300270000",
    1009 => x"000bff9c00240000",
    1010 => x"fff5ff9c00240000",
    1011 => x"fff5ffa300270000",
    1012 => x"fff5ffa300270000",
    1013 => x"fff5ffa4002e0000",
    1014 => x"0000ffa0002d0000",
    1015 => x"0000ff9f00260000",
    1016 => x"0000ff9f00260000",
    1017 => x"000bffa300270000",
    1018 => x"fff5ffa300270000",
    1019 => x"0000ff9f00260000",
    1020 => x"0000ff9f00260000",
    1021 => x"0000ff9700230000",
    1022 => x"0005ff9700230000",
    1023 => x"000bffa300270000",
    1024 => x"fff5ffa300270000",
    1025 => x"fffbff9700230000",
    1026 => x"0014001100340000",
    1027 => x"000f001000310000",
    1028 => x"0013000800300000",
    1029 => x"0015000a00330000",
    1030 => x"0015000a00330000",
    1031 => x"0014001100340000",
    1032 => x"ffec001100340000",
    1033 => x"ffeb000a00330000",
    1034 => x"ffeb000a00330000",
    1035 => x"ffed000800300000",
    1036 => x"fff1001000310000",
    1037 => x"ffec001100340000",
    1038 => x"0014001a00340000",
    1039 => x"000e001b00320000",
    1040 => x"0014001100340000",
    1041 => x"0014001a00340000",
    1042 => x"ffec001a00340000",
    1043 => x"ffec001100340000",
    1044 => x"fff2001b00320000",
    1045 => x"ffec001a00340000",
    1046 => x"0018002300340000",
    1047 => x"0013002700330000",
    1048 => x"0014001a00340000",
    1049 => x"0018002300340000",
    1050 => x"ffe8002300340000",
    1051 => x"ffec001a00340000",
    1052 => x"ffed002700330000",
    1053 => x"ffe8002300340000",
    1054 => x"0017000300300000",
    1055 => x"001a000500340000",
    1056 => x"001a000500340000",
    1057 => x"0015000a00330000",
    1058 => x"ffeb000a00330000",
    1059 => x"ffe6000500340000",
    1060 => x"ffe6000500340000",
    1061 => x"ffe9000300300000",
    1062 => x"002bfffa002b0000",
    1063 => x"002bffff00300000",
    1064 => x"002bffff00300000",
    1065 => x"001a000500340000",
    1066 => x"ffe6000500340000",
    1067 => x"ffd5ffff00300000",
    1068 => x"ffd5ffff00300000",
    1069 => x"ffd5fffa002b0000",
    1070 => x"0038ffff00280000",
    1071 => x"00360004002d0000",
    1072 => x"00360004002d0000",
    1073 => x"002bffff00300000",
    1074 => x"ffd5ffff00300000",
    1075 => x"ffca0004002d0000",
    1076 => x"ffca0004002d0000",
    1077 => x"ffc8ffff00280000",
    1078 => x"0047000e00250000",
    1079 => x"0042000f00280000",
    1080 => x"0042000f00280000",
    1081 => x"00360004002d0000",
    1082 => x"ffca0004002d0000",
    1083 => x"ffbe000f00280000",
    1084 => x"ffbe000f00280000",
    1085 => x"ffb9000e00250000",
    1086 => x"0049001a00250000",
    1087 => x"0043001900290000",
    1088 => x"0043001900290000",
    1089 => x"0042000f00280000",
    1090 => x"ffbe000f00280000",
    1091 => x"ffbd001900290000",
    1092 => x"ffbd001900290000",
    1093 => x"ffb7001a00250000",
    1094 => x"0044002300270000",
    1095 => x"00400020002a0000",
    1096 => x"00400020002a0000",
    1097 => x"0043001900290000",
    1098 => x"ffbd001900290000",
    1099 => x"ffc00020002a0000",
    1100 => x"ffc00020002a0000",
    1101 => x"ffbc002300270000",
    1102 => x"0031002a002d0000",
    1103 => x"0030002600330000",
    1104 => x"0030002600330000",
    1105 => x"00400020002a0000",
    1106 => x"ffc00020002a0000",
    1107 => x"ffd0002600330000",
    1108 => x"ffd0002600330000",
    1109 => x"ffcf002a002d0000",
    1110 => x"0025002f00300000",
    1111 => x"0026002900310000",
    1112 => x"0026002900310000",
    1113 => x"0030002600330000",
    1114 => x"ffd0002600330000",
    1115 => x"ffda002900310000",
    1116 => x"ffda002900310000",
    1117 => x"ffdb002f00300000",
    1118 => x"001c002e00310000",
    1119 => x"001f002800330000",
    1120 => x"001f002800330000",
    1121 => x"0026002900310000",
    1122 => x"ffda002900310000",
    1123 => x"ffe1002800330000",
    1124 => x"ffe1002800330000",
    1125 => x"ffe4002e00310000",
    1126 => x"0018002300340000",
    1127 => x"001f002800330000",
    1128 => x"ffe1002800330000",
    1129 => x"ffe8002300340000",
    1130 => x"0020002600320000",
    1131 => x"001f002800330000",
    1132 => x"0018002300340000",
    1133 => x"001b002100310000",
    1134 => x"001b002100310000",
    1135 => x"0020002600320000",
    1136 => x"ffe0002600320000",
    1137 => x"ffe5002100310000",
    1138 => x"ffe5002100310000",
    1139 => x"ffe8002300340000",
    1140 => x"ffe1002800330000",
    1141 => x"ffe0002600320000",
    1142 => x"0026002700300000",
    1143 => x"0026002900310000",
    1144 => x"0020002600320000",
    1145 => x"0026002700300000",
    1146 => x"ffda002700300000",
    1147 => x"ffe0002600320000",
    1148 => x"ffda002900310000",
    1149 => x"ffda002700300000",
    1150 => x"002f002500300000",
    1151 => x"0030002600330000",
    1152 => x"0026002700300000",
    1153 => x"002f002500300000",
    1154 => x"ffd1002500300000",
    1155 => x"ffda002700300000",
    1156 => x"ffd0002600330000",
    1157 => x"ffd1002500300000",
    1158 => x"003c001f00280000",
    1159 => x"00400020002a0000",
    1160 => x"002f002500300000",
    1161 => x"003c001f00280000",
    1162 => x"ffc4001f00280000",
    1163 => x"ffd1002500300000",
    1164 => x"ffc00020002a0000",
    1165 => x"ffc4001f00280000",
    1166 => x"003f001800280000",
    1167 => x"0043001900290000",
    1168 => x"003c001f00280000",
    1169 => x"003f001800280000",
    1170 => x"ffc1001800280000",
    1171 => x"ffc4001f00280000",
    1172 => x"ffbd001900290000",
    1173 => x"ffc1001800280000",
    1174 => x"003e001000280000",
    1175 => x"0042000f00280000",
    1176 => x"003f001800280000",
    1177 => x"003e001000280000",
    1178 => x"ffc2001000280000",
    1179 => x"ffc1001800280000",
    1180 => x"ffbe000f00280000",
    1181 => x"ffc2001000280000",
    1182 => x"00340006002b0000",
    1183 => x"00360004002d0000",
    1184 => x"003e001000280000",
    1185 => x"00340006002b0000",
    1186 => x"ffcc0006002b0000",
    1187 => x"ffc2001000280000",
    1188 => x"ffca0004002d0000",
    1189 => x"ffcc0006002b0000",
    1190 => x"002b0002002e0000",
    1191 => x"002bffff00300000",
    1192 => x"00340006002b0000",
    1193 => x"002b0002002e0000",
    1194 => x"ffd50002002e0000",
    1195 => x"ffcc0006002b0000",
    1196 => x"ffd5ffff00300000",
    1197 => x"ffd50002002e0000",
    1198 => x"001c000700310000",
    1199 => x"001a000500340000",
    1200 => x"002b0002002e0000",
    1201 => x"001c000700310000",
    1202 => x"ffe4000700310000",
    1203 => x"ffd50002002e0000",
    1204 => x"ffe6000500340000",
    1205 => x"ffe4000700310000",
    1206 => x"0017000c00300000",
    1207 => x"0015000a00330000",
    1208 => x"001c000700310000",
    1209 => x"0017000c00300000",
    1210 => x"ffe9000c00300000",
    1211 => x"ffe4000700310000",
    1212 => x"ffeb000a00330000",
    1213 => x"ffe9000c00300000",
    1214 => x"0014001a00340000",
    1215 => x"0016001a00310000",
    1216 => x"0016001a00310000",
    1217 => x"001b002100310000",
    1218 => x"ffe5002100310000",
    1219 => x"ffea001a00310000",
    1220 => x"ffea001a00310000",
    1221 => x"ffec001a00340000",
    1222 => x"0014001100340000",
    1223 => x"0016001200300000",
    1224 => x"0016001200300000",
    1225 => x"0016001a00310000",
    1226 => x"ffea001a00310000",
    1227 => x"ffea001200300000",
    1228 => x"ffea001200300000",
    1229 => x"ffec001100340000",
    1230 => x"0017000c00300000",
    1231 => x"0016001200300000",
    1232 => x"ffea001200300000",
    1233 => x"ffe9000c00300000",
    1234 => x"0000002700200000",
    1235 => x"0000002900300000",
    1236 => x"0007003000300000",
    1237 => x"000c002d00200000",
    1238 => x"000c002d00200000",
    1239 => x"0000002700200000",
    1240 => x"0000002700200000",
    1241 => x"fff4002d00200000",
    1242 => x"fff4002d00200000",
    1243 => x"fff9003000300000",
    1244 => x"0012004a00310000",
    1245 => x"0016004400210000",
    1246 => x"0016004400210000",
    1247 => x"000c002d00200000",
    1248 => x"fff4002d00200000",
    1249 => x"ffea004400210000",
    1250 => x"ffea004400210000",
    1251 => x"ffee004a00310000",
    1252 => x"0024004e002f0000",
    1253 => x"00260047001f0000",
    1254 => x"00260047001f0000",
    1255 => x"0016004400210000",
    1256 => x"ffea004400210000",
    1257 => x"ffda0047001f0000",
    1258 => x"ffda0047001f0000",
    1259 => x"ffdc004e002f0000",
    1260 => x"0038003d00290000",
    1261 => x"00370037001a0000",
    1262 => x"00370037001a0000",
    1263 => x"00260047001f0000",
    1264 => x"ffda0047001f0000",
    1265 => x"ffc90037001a0000",
    1266 => x"ffc90037001a0000",
    1267 => x"ffc8003d00290000",
    1268 => x"0051002f00220000",
    1269 => x"004d002c00130000",
    1270 => x"004d002c00130000",
    1271 => x"00370037001a0000",
    1272 => x"ffc90037001a0000",
    1273 => x"ffb3002c00130000",
    1274 => x"ffb3002c00130000",
    1275 => x"ffaf002f00220000",
    1276 => x"00620029001f0000",
    1277 => x"005b002700100000",
    1278 => x"005b002700100000",
    1279 => x"004d002c00130000",
    1280 => x"ffb3002c00130000",
    1281 => x"ffa5002700100000",
    1282 => x"ffa5002700100000",
    1283 => x"ff9e0029001f0000",
    1284 => x"005e0009000e0000",
    1285 => x"0058000b00060000",
    1286 => x"0058000b00060000",
    1287 => x"005b002700100000",
    1288 => x"ffa5002700100000",
    1289 => x"ffa8000b00060000",
    1290 => x"ffa8000b00060000",
    1291 => x"ffa20009000e0000",
    1292 => x"0048fff400180000",
    1293 => x"0044fff8000a0000",
    1294 => x"0044fff8000a0000",
    1295 => x"0058000b00060000",
    1296 => x"ffa8000b00060000",
    1297 => x"ffbcfff8000a0000",
    1298 => x"ffbcfff8000a0000",
    1299 => x"ffb8fff400180000",
    1300 => x"0032ffe800180000",
    1301 => x"0032ffee00100000",
    1302 => x"0032ffee00100000",
    1303 => x"0044fff8000a0000",
    1304 => x"ffbcfff8000a0000",
    1305 => x"ffceffee00100000",
    1306 => x"ffceffee00100000",
    1307 => x"ffceffe800180000",
    1308 => x"000effbb00040000",
    1309 => x"0000ffb700000000",
    1310 => x"0000ffb700000000",
    1311 => x"0000ffc1fffb0000",
    1312 => x"0000ffc1fffb0000",
    1313 => x"0014ffc9fff90000",
    1314 => x"0014ffc9fff90000",
    1315 => x"000effbb00040000",
    1316 => x"fff2ffbb00040000",
    1317 => x"ffecffc9fff90000",
    1318 => x"ffecffc9fff90000",
    1319 => x"0000ffc1fffb0000",
    1320 => x"0000ffb700000000",
    1321 => x"fff2ffbb00040000",
    1322 => x"0010ffa200050000",
    1323 => x"0000ff9d00020000",
    1324 => x"0000ff9d00020000",
    1325 => x"0000ffb700000000",
    1326 => x"000effbb00040000",
    1327 => x"0010ffa200050000",
    1328 => x"fff0ffa200050000",
    1329 => x"fff2ffbb00040000",
    1330 => x"0000ff9d00020000",
    1331 => x"fff0ffa200050000",
    1332 => x"0013ff8d000d0000",
    1333 => x"0000ff8900100000",
    1334 => x"0000ff8900100000",
    1335 => x"0000ff9d00020000",
    1336 => x"0010ffa200050000",
    1337 => x"0013ff8d000d0000",
    1338 => x"ffedff8d000d0000",
    1339 => x"fff0ffa200050000",
    1340 => x"0000ff8900100000",
    1341 => x"ffedff8d000d0000",
    1342 => x"0013ff8d000d0000",
    1343 => x"0014ff8a001a0000",
    1344 => x"0000ff88001d0000",
    1345 => x"0000ff8900100000",
    1346 => x"ffecff8a001a0000",
    1347 => x"ffedff8d000d0000",
    1348 => x"0025ff9000080000",
    1349 => x"0025ff8d00170000",
    1350 => x"0013ff8d000d0000",
    1351 => x"0025ff9000080000",
    1352 => x"ffdbff9000080000",
    1353 => x"ffedff8d000d0000",
    1354 => x"ffdbff8d00170000",
    1355 => x"ffdbff9000080000",
    1356 => x"0021ffa700070000",
    1357 => x"002aff9300180000",
    1358 => x"0025ff9000080000",
    1359 => x"0021ffa700070000",
    1360 => x"ffdfffa700070000",
    1361 => x"ffdbff9000080000",
    1362 => x"ffd6ff9300180000",
    1363 => x"ffdfffa700070000",
    1364 => x"001cffbf00080000",
    1365 => x"0028ffa9001c0000",
    1366 => x"0021ffa700070000",
    1367 => x"001cffbf00080000",
    1368 => x"ffe4ffbf00080000",
    1369 => x"ffdfffa700070000",
    1370 => x"ffd8ffa9001c0000",
    1371 => x"ffe4ffbf00080000",
    1372 => x"0021ffa700070000",
    1373 => x"0010ffa200050000",
    1374 => x"000effbb00040000",
    1375 => x"001cffbf00080000",
    1376 => x"ffe4ffbf00080000",
    1377 => x"fff2ffbb00040000",
    1378 => x"fff0ffa200050000",
    1379 => x"ffdfffa700070000",
    1380 => x"0014ffc9fff90000",
    1381 => x"001bffd000090000",
    1382 => x"001bffd000090000",
    1383 => x"001cffbf00080000",
    1384 => x"ffe4ffbf00080000",
    1385 => x"ffe5ffd000090000",
    1386 => x"ffe5ffd000090000",
    1387 => x"ffecffc9fff90000",
    1388 => x"001bffd000090000",
    1389 => x"0024ffc7001c0000",
    1390 => x"ffdcffc7001c0000",
    1391 => x"ffe5ffd000090000",
    1392 => x"001dffd5001a0000",
    1393 => x"0019ffd8000c0000",
    1394 => x"0019ffd8000c0000",
    1395 => x"0018ffdf00100000",
    1396 => x"0018ffdf00100000",
    1397 => x"001bffdc001a0000",
    1398 => x"ffe5ffdc001a0000",
    1399 => x"ffe8ffdf00100000",
    1400 => x"ffe8ffdf00100000",
    1401 => x"ffe7ffd8000c0000",
    1402 => x"ffe7ffd8000c0000",
    1403 => x"ffe3ffd5001a0000",
    1404 => x"001bffd000090000",
    1405 => x"0019ffd8000c0000",
    1406 => x"ffe7ffd8000c0000",
    1407 => x"ffe5ffd000090000",
    1408 => x"0017ffe500140000",
    1409 => x"0017ffe3001b0000",
    1410 => x"0018ffdf00100000",
    1411 => x"0017ffe500140000",
    1412 => x"ffe9ffe500140000",
    1413 => x"ffe8ffdf00100000",
    1414 => x"ffe9ffe3001b0000",
    1415 => x"ffe9ffe500140000",
    1416 => x"0017ffe500140000",
    1417 => x"0032ffee00100000",
    1418 => x"ffceffee00100000",
    1419 => x"ffe9ffe500140000",
    1420 => x"0000ffe2ff8f0000",
    1421 => x"00000000ff7d0000",
    1422 => x"00000000ff7d0000",
    1423 => x"0026ffffff900000",
    1424 => x"0026ffffff900000",
    1425 => x"0027ffe7ff9e0000",
    1426 => x"0027ffe7ff9e0000",
    1427 => x"0000ffe2ff8f0000",
    1428 => x"0000ffe2ff8f0000",
    1429 => x"ffd9ffe7ff9e0000",
    1430 => x"ffd9ffe7ff9e0000",
    1431 => x"ffdaffffff900000",
    1432 => x"ffdaffffff900000",
    1433 => x"00000000ff7d0000",
    1434 => x"0000ffcdffb30000",
    1435 => x"0000ffe2ff8f0000",
    1436 => x"0027ffe7ff9e0000",
    1437 => x"0022ffd5ffbd0000",
    1438 => x"0022ffd5ffbd0000",
    1439 => x"0000ffcdffb30000",
    1440 => x"0000ffcdffb30000",
    1441 => x"ffdeffd5ffbd0000",
    1442 => x"ffdeffd5ffbd0000",
    1443 => x"ffd9ffe7ff9e0000",
    1444 => x"0000ffc4fff10000",
    1445 => x"0000ffcdffb30000",
    1446 => x"0022ffd5ffbd0000",
    1447 => x"0018ffccffee0000",
    1448 => x"0018ffccffee0000",
    1449 => x"0000ffc4fff10000",
    1450 => x"0000ffc4fff10000",
    1451 => x"ffe8ffccffee0000",
    1452 => x"ffe8ffccffee0000",
    1453 => x"ffdeffd5ffbd0000",
    1454 => x"0000ffc1fffb0000",
    1455 => x"0000ffc4fff10000",
    1456 => x"0018ffccffee0000",
    1457 => x"0014ffc9fff90000",
    1458 => x"ffecffc9fff90000",
    1459 => x"ffe8ffccffee0000",
    1460 => x"0018ffccffee0000",
    1461 => x"0019ffd8000c0000",
    1462 => x"ffe7ffd8000c0000",
    1463 => x"ffe8ffccffee0000",
    1464 => x"00610013ffe10000",
    1465 => x"0058000b00060000",
    1466 => x"0044fff8000a0000",
    1467 => x"0054fff3ffe30000",
    1468 => x"0054fff3ffe30000",
    1469 => x"00610013ffe10000",
    1470 => x"ff9f0013ffe10000",
    1471 => x"ffacfff3ffe30000",
    1472 => x"ffacfff3ffe30000",
    1473 => x"ffbcfff8000a0000",
    1474 => x"ffa8000b00060000",
    1475 => x"ff9f0013ffe10000",
    1476 => x"00000000ff7d0000",
    1477 => x"00000038ff7a0000",
    1478 => x"00000038ff7a0000",
    1479 => x"0034002aff8b0000",
    1480 => x"0034002aff8b0000",
    1481 => x"0026ffffff900000",
    1482 => x"ffdaffffff900000",
    1483 => x"ffcc002aff8b0000",
    1484 => x"ffcc002aff8b0000",
    1485 => x"00000038ff7a0000",
    1486 => x"00000068ffd20000",
    1487 => x"0000005efffc0000",
    1488 => x"0000005efffc0000",
    1489 => x"00340059fff60000",
    1490 => x"00340059fff60000",
    1491 => x"00340062ffd30000",
    1492 => x"00340062ffd30000",
    1493 => x"00000068ffd20000",
    1494 => x"00000068ffd20000",
    1495 => x"ffcc0062ffd30000",
    1496 => x"ffcc0062ffd30000",
    1497 => x"ffcc0059fff60000",
    1498 => x"ffcc0059fff60000",
    1499 => x"0000005efffc0000",
    1500 => x"0000005eff9d0000",
    1501 => x"00000068ffd20000",
    1502 => x"00340062ffd30000",
    1503 => x"0034005bffb00000",
    1504 => x"0034005bffb00000",
    1505 => x"0000005eff9d0000",
    1506 => x"0000005eff9d0000",
    1507 => x"ffcc005bffb00000",
    1508 => x"ffcc005bffb00000",
    1509 => x"ffcc0062ffd30000",
    1510 => x"00000038ff7a0000",
    1511 => x"0000005eff9d0000",
    1512 => x"0034005bffb00000",
    1513 => x"0034002aff8b0000",
    1514 => x"ffcc002aff8b0000",
    1515 => x"ffcc005bffb00000",
    1516 => x"0048002cfffb0000",
    1517 => x"004d002c00130000",
    1518 => x"005b002700100000",
    1519 => x"0053002700010000",
    1520 => x"0053002700010000",
    1521 => x"0048002cfffb0000",
    1522 => x"ffb8002cfffb0000",
    1523 => x"ffad002700010000",
    1524 => x"ffad002700010000",
    1525 => x"ffa5002700100000",
    1526 => x"ffb3002c00130000",
    1527 => x"ffb8002cfffb0000",
    1528 => x"00490048ffe10000",
    1529 => x"0048002cfffb0000",
    1530 => x"0053002700010000",
    1531 => x"005b0038ffe90000",
    1532 => x"005b0038ffe90000",
    1533 => x"00490048ffe10000",
    1534 => x"ffb70048ffe10000",
    1535 => x"ffa50038ffe90000",
    1536 => x"ffa50038ffe90000",
    1537 => x"ffad002700010000",
    1538 => x"ffb8002cfffb0000",
    1539 => x"ffb70048ffe10000",
    1540 => x"0049004effc50000",
    1541 => x"00490048ffe10000",
    1542 => x"005b0038ffe90000",
    1543 => x"005b003fffce0000",
    1544 => x"005b003fffce0000",
    1545 => x"0049004effc50000",
    1546 => x"ffb7004effc50000",
    1547 => x"ffa5003fffce0000",
    1548 => x"ffa5003fffce0000",
    1549 => x"ffa50038ffe90000",
    1550 => x"ffb70048ffe10000",
    1551 => x"ffb7004effc50000",
    1552 => x"00490046ffa90000",
    1553 => x"0049004effc50000",
    1554 => x"005b003fffce0000",
    1555 => x"005b0036ffb20000",
    1556 => x"005b0036ffb20000",
    1557 => x"00490046ffa90000",
    1558 => x"ffb70046ffa90000",
    1559 => x"ffa50036ffb20000",
    1560 => x"ffa50036ffb20000",
    1561 => x"ffa5003fffce0000",
    1562 => x"ffb7004effc50000",
    1563 => x"ffb70046ffa90000",
    1564 => x"005b0036ffb20000",
    1565 => x"00580017ffa90000",
    1566 => x"00580017ffa90000",
    1567 => x"0046001eff990000",
    1568 => x"0046001eff990000",
    1569 => x"00490046ffa90000",
    1570 => x"ffb70046ffa90000",
    1571 => x"ffba001eff990000",
    1572 => x"ffba001eff990000",
    1573 => x"ffa80017ffa90000",
    1574 => x"ffa80017ffa90000",
    1575 => x"ffa50036ffb20000",
    1576 => x"0046001eff990000",
    1577 => x"0034002aff8b0000",
    1578 => x"0034005bffb00000",
    1579 => x"00490046ffa90000",
    1580 => x"ffb70046ffa90000",
    1581 => x"ffcc005bffb00000",
    1582 => x"ffcc002aff8b0000",
    1583 => x"ffba001eff990000",
    1584 => x"00340062ffd30000",
    1585 => x"0049004effc50000",
    1586 => x"ffb7004effc50000",
    1587 => x"ffcc0062ffd30000",
    1588 => x"00340059fff60000",
    1589 => x"00490048ffe10000",
    1590 => x"ffb70048ffe10000",
    1591 => x"ffcc0059fff60000",
    1592 => x"00340059fff60000",
    1593 => x"00340034000c0000",
    1594 => x"00340034000c0000",
    1595 => x"0048002cfffb0000",
    1596 => x"ffb8002cfffb0000",
    1597 => x"ffcc0034000c0000",
    1598 => x"ffcc0034000c0000",
    1599 => x"ffcc0059fff60000",
    1600 => x"00340034000c0000",
    1601 => x"00370037001a0000",
    1602 => x"ffc90037001a0000",
    1603 => x"ffcc0034000c0000",
    1604 => x"0000005efffc0000",
    1605 => x"00000039001c0000",
    1606 => x"00000039001c0000",
    1607 => x"00340034000c0000",
    1608 => x"ffcc0034000c0000",
    1609 => x"00000039001c0000",
    1610 => x"00370037001a0000",
    1611 => x"000c002d00200000",
    1612 => x"fff4002d00200000",
    1613 => x"ffc90037001a0000",
    1614 => x"00000039001c0000",
    1615 => x"000c002d00200000",
    1616 => x"fff4002d00200000",
    1617 => x"00000039001c0000",
    1618 => x"00000039001c0000",
    1619 => x"0000002700200000",
    1620 => x"00610013ffe10000",
    1621 => x"0053002700010000",
    1622 => x"ffad002700010000",
    1623 => x"ff9f0013ffe10000",
    1624 => x"00610013ffe10000",
    1625 => x"0062001dffd60000",
    1626 => x"0062001dffd60000",
    1627 => x"005b0038ffe90000",
    1628 => x"ffa50038ffe90000",
    1629 => x"ff9e001dffd60000",
    1630 => x"ff9e001dffd60000",
    1631 => x"ff9f0013ffe10000",
    1632 => x"0062001dffd60000",
    1633 => x"005d001effc40000",
    1634 => x"005d001effc40000",
    1635 => x"005b003fffce0000",
    1636 => x"ffa5003fffce0000",
    1637 => x"ffa3001effc40000",
    1638 => x"ffa3001effc40000",
    1639 => x"ff9e001dffd60000",
    1640 => x"005d001effc40000",
    1641 => x"00580017ffa90000",
    1642 => x"ffa80017ffa90000",
    1643 => x"ffa3001effc40000",
    1644 => x"002effe5ffec0000",
    1645 => x"0018ffccffee0000",
    1646 => x"0022ffd5ffbd0000",
    1647 => x"0031ffe2ffc30000",
    1648 => x"0031ffe2ffc30000",
    1649 => x"002effe5ffec0000",
    1650 => x"ffd2ffe5ffec0000",
    1651 => x"ffcfffe2ffc30000",
    1652 => x"ffcfffe2ffc30000",
    1653 => x"ffdeffd5ffbd0000",
    1654 => x"ffe8ffccffee0000",
    1655 => x"ffd2ffe5ffec0000",
    1656 => x"0044ffeaffc90000",
    1657 => x"0054fff3ffe30000",
    1658 => x"0054fff3ffe30000",
    1659 => x"002effe5ffec0000",
    1660 => x"0031ffe2ffc30000",
    1661 => x"0044ffeaffc90000",
    1662 => x"ffbcffeaffc90000",
    1663 => x"ffcfffe2ffc30000",
    1664 => x"ffd2ffe5ffec0000",
    1665 => x"ffacfff3ffe30000",
    1666 => x"ffacfff3ffe30000",
    1667 => x"ffbcffeaffc90000",
    1668 => x"0032ffee00100000",
    1669 => x"002effe5ffec0000",
    1670 => x"ffd2ffe5ffec0000",
    1671 => x"ffceffee00100000",
    1672 => x"0032ffee00100000",
    1673 => x"0018ffdf00100000",
    1674 => x"0019ffd8000c0000",
    1675 => x"002effe5ffec0000",
    1676 => x"ffd2ffe5ffec0000",
    1677 => x"ffe7ffd8000c0000",
    1678 => x"ffe8ffdf00100000",
    1679 => x"ffceffee00100000",
    1680 => x"00580017ffa90000",
    1681 => x"0049fff7ffaa0000",
    1682 => x"0049fff7ffaa0000",
    1683 => x"0037fffbff9d0000",
    1684 => x"0037fffbff9d0000",
    1685 => x"0046001eff990000",
    1686 => x"ffba001eff990000",
    1687 => x"ffc9fffbff9d0000",
    1688 => x"ffc9fffbff9d0000",
    1689 => x"ffb7fff7ffaa0000",
    1690 => x"ffb7fff7ffaa0000",
    1691 => x"ffa80017ffa90000",
    1692 => x"0037fffbff9d0000",
    1693 => x"0026ffffff900000",
    1694 => x"ffdaffffff900000",
    1695 => x"ffc9fffbff9d0000",
    1696 => x"0049fff7ffaa0000",
    1697 => x"0044ffeaffc90000",
    1698 => x"0031ffe2ffc30000",
    1699 => x"0037fffbff9d0000",
    1700 => x"ffc9fffbff9d0000",
    1701 => x"ffcfffe2ffc30000",
    1702 => x"ffbcffeaffc90000",
    1703 => x"ffb7fff7ffaa0000",
    1704 => x"0027ffe7ff9e0000",
    1705 => x"0037fffbff9d0000",
    1706 => x"ffc9fffbff9d0000",
    1707 => x"ffd9ffe7ff9e0000",
    1708 => x"00730027ffba0000",
    1709 => x"0074002fffb80000",
    1710 => x"0074002fffb80000",
    1711 => x"00650027ffc10000",
    1712 => x"00650027ffc10000",
    1713 => x"00690021ffc20000",
    1714 => x"00690021ffc20000",
    1715 => x"00730027ffba0000",
    1716 => x"ff8d0027ffba0000",
    1717 => x"ff970021ffc20000",
    1718 => x"ff970021ffc20000",
    1719 => x"ff9b0027ffc10000",
    1720 => x"ff9b0027ffc10000",
    1721 => x"ff8c002fffb80000",
    1722 => x"ff8c002fffb80000",
    1723 => x"ff8d0027ffba0000",
    1724 => x"008c0032ffab0000",
    1725 => x"0074002fffb80000",
    1726 => x"00730027ffba0000",
    1727 => x"0087002affaf0000",
    1728 => x"0087002affaf0000",
    1729 => x"008c0032ffab0000",
    1730 => x"ff740032ffab0000",
    1731 => x"ff79002affaf0000",
    1732 => x"ff79002affaf0000",
    1733 => x"ff8d0027ffba0000",
    1734 => x"ff8c002fffb80000",
    1735 => x"ff740032ffab0000",
    1736 => x"009a001dffab0000",
    1737 => x"008c0032ffab0000",
    1738 => x"0087002affaf0000",
    1739 => x"00900019ffad0000",
    1740 => x"00900019ffad0000",
    1741 => x"009a001dffab0000",
    1742 => x"ff66001dffab0000",
    1743 => x"ff700019ffad0000",
    1744 => x"ff700019ffad0000",
    1745 => x"ff79002affaf0000",
    1746 => x"ff740032ffab0000",
    1747 => x"ff66001dffab0000",
    1748 => x"0092ffffffaa0000",
    1749 => x"009a001dffab0000",
    1750 => x"00900019ffad0000",
    1751 => x"008a0001ffad0000",
    1752 => x"008a0001ffad0000",
    1753 => x"0092ffffffaa0000",
    1754 => x"ff6effffffaa0000",
    1755 => x"ff760001ffad0000",
    1756 => x"ff760001ffad0000",
    1757 => x"ff700019ffad0000",
    1758 => x"ff66001dffab0000",
    1759 => x"ff6effffffaa0000",
    1760 => x"0076ffedffb60000",
    1761 => x"0092ffffffaa0000",
    1762 => x"008a0001ffad0000",
    1763 => x"0075fff4ffb90000",
    1764 => x"0075fff4ffb90000",
    1765 => x"0076ffedffb60000",
    1766 => x"ff8affedffb60000",
    1767 => x"ff8bfff4ffb90000",
    1768 => x"ff8bfff4ffb90000",
    1769 => x"ff760001ffad0000",
    1770 => x"ff6effffffaa0000",
    1771 => x"ff8affedffb60000",
    1772 => x"0058ffe8ffcd0000",
    1773 => x"0076ffedffb60000",
    1774 => x"0075fff4ffb90000",
    1775 => x"005efff0ffcc0000",
    1776 => x"005efff0ffcc0000",
    1777 => x"0058ffe8ffcd0000",
    1778 => x"ffa8ffe8ffcd0000",
    1779 => x"ffa2fff0ffcc0000",
    1780 => x"ffa2fff0ffcc0000",
    1781 => x"ff8bfff4ffb90000",
    1782 => x"ff8affedffb60000",
    1783 => x"ffa8ffe8ffcd0000",
    1784 => x"0075fff4ffb90000",
    1785 => x"0076fff8ffb10000",
    1786 => x"0076fff8ffb10000",
    1787 => x"0064fff6ffc30000",
    1788 => x"0064fff6ffc30000",
    1789 => x"005efff0ffcc0000",
    1790 => x"ffa2fff0ffcc0000",
    1791 => x"ff9cfff6ffc30000",
    1792 => x"ff9cfff6ffc30000",
    1793 => x"ff8afff8ffb10000",
    1794 => x"ff8afff8ffb10000",
    1795 => x"ff8bfff4ffb90000",
    1796 => x"008a0001ffad0000",
    1797 => x"00870003ffa90000",
    1798 => x"00870003ffa90000",
    1799 => x"0076fff8ffb10000",
    1800 => x"ff8afff8ffb10000",
    1801 => x"ff790003ffa90000",
    1802 => x"ff790003ffa90000",
    1803 => x"ff760001ffad0000",
    1804 => x"00900019ffad0000",
    1805 => x"008c0015ffa90000",
    1806 => x"008c0015ffa90000",
    1807 => x"00870003ffa90000",
    1808 => x"ff790003ffa90000",
    1809 => x"ff740015ffa90000",
    1810 => x"ff740015ffa90000",
    1811 => x"ff700019ffad0000",
    1812 => x"0087002affaf0000",
    1813 => x"00850021ffa90000",
    1814 => x"00850021ffa90000",
    1815 => x"008c0015ffa90000",
    1816 => x"ff740015ffa90000",
    1817 => x"ff7b0021ffa90000",
    1818 => x"ff7b0021ffa90000",
    1819 => x"ff79002affaf0000",
    1820 => x"00730027ffba0000",
    1821 => x"0074001fffb20000",
    1822 => x"0074001fffb20000",
    1823 => x"00850021ffa90000",
    1824 => x"ff7b0021ffa90000",
    1825 => x"ff8c001fffb20000",
    1826 => x"ff8c001fffb20000",
    1827 => x"ff8d0027ffba0000",
    1828 => x"00690021ffc20000",
    1829 => x"006b001bffba0000",
    1830 => x"006b001bffba0000",
    1831 => x"0074001fffb20000",
    1832 => x"ff8c001fffb20000",
    1833 => x"ff95001bffba0000",
    1834 => x"ff95001bffba0000",
    1835 => x"ff970021ffc20000",
    1836 => x"0053fff8ffd30000",
    1837 => x"0054fff3ffe30000",
    1838 => x"0044ffeaffc90000",
    1839 => x"0052fff6ffc80000",
    1840 => x"0052fff6ffc80000",
    1841 => x"0053fff8ffd30000",
    1842 => x"ffadfff8ffd30000",
    1843 => x"ffaefff6ffc80000",
    1844 => x"ffaefff6ffc80000",
    1845 => x"ffbcffeaffc90000",
    1846 => x"ffacfff3ffe30000",
    1847 => x"ffadfff8ffd30000",
    1848 => x"0044ffeaffc90000",
    1849 => x"0058ffe8ffcd0000",
    1850 => x"005efff0ffcc0000",
    1851 => x"0052fff6ffc80000",
    1852 => x"ffaefff6ffc80000",
    1853 => x"ffa2fff0ffcc0000",
    1854 => x"ffa8ffe8ffcd0000",
    1855 => x"ffbcffeaffc90000",
    1856 => x"0053fff8ffd30000",
    1857 => x"0062001dffd60000",
    1858 => x"ff9e001dffd60000",
    1859 => x"ffadfff8ffd30000",
    1860 => x"00650027ffc10000",
    1861 => x"005d001effc40000",
    1862 => x"005d001effc40000",
    1863 => x"00600019ffc30000",
    1864 => x"00600019ffc30000",
    1865 => x"00690021ffc20000",
    1866 => x"ff970021ffc20000",
    1867 => x"ffa00019ffc30000",
    1868 => x"ffa00019ffc30000",
    1869 => x"ffa3001effc40000",
    1870 => x"ffa3001effc40000",
    1871 => x"ff9b0027ffc10000",
    1872 => x"0064fff6ffc30000",
    1873 => x"005cfff7ffbc0000",
    1874 => x"005cfff7ffbc0000",
    1875 => x"0052fff6ffc80000",
    1876 => x"ffaefff6ffc80000",
    1877 => x"ffa4fff7ffbc0000",
    1878 => x"ffa4fff7ffbc0000",
    1879 => x"ff9cfff6ffc30000",
    1880 => x"005cfff7ffbc0000",
    1881 => x"0060fffaffbc0000",
    1882 => x"0060fffaffbc0000",
    1883 => x"0052fffdffc60000",
    1884 => x"0052fffdffc60000",
    1885 => x"0052fff6ffc80000",
    1886 => x"ffaefff6ffc80000",
    1887 => x"ffaefffdffc60000",
    1888 => x"ffaefffdffc60000",
    1889 => x"ffa0fffaffbc0000",
    1890 => x"ffa0fffaffbc0000",
    1891 => x"ffa4fff7ffbc0000",
    1892 => x"005d0002ffbc0000",
    1893 => x"00560003ffbc0000",
    1894 => x"00560003ffbc0000",
    1895 => x"0052fffdffc60000",
    1896 => x"0060fffaffbc0000",
    1897 => x"005d0002ffbc0000",
    1898 => x"ffa30002ffbc0000",
    1899 => x"ffa0fffaffbc0000",
    1900 => x"ffaefffdffc60000",
    1901 => x"ffaa0003ffbc0000",
    1902 => x"ffaa0003ffbc0000",
    1903 => x"ffa30002ffbc0000",
    1904 => x"00560003ffbc0000",
    1905 => x"005f000cffbc0000",
    1906 => x"005f000cffbc0000",
    1907 => x"005b000fffc30000",
    1908 => x"005b000fffc30000",
    1909 => x"0052fffdffc60000",
    1910 => x"ffaefffdffc60000",
    1911 => x"ffa5000fffc30000",
    1912 => x"ffa5000fffc30000",
    1913 => x"ffa1000cffbc0000",
    1914 => x"ffa1000cffbc0000",
    1915 => x"ffaa0003ffbc0000",
    1916 => x"00650014ffbd0000",
    1917 => x"00600019ffc30000",
    1918 => x"00600019ffc30000",
    1919 => x"005b000fffc30000",
    1920 => x"005f000cffbc0000",
    1921 => x"00650014ffbd0000",
    1922 => x"ff9b0014ffbd0000",
    1923 => x"ffa1000cffbc0000",
    1924 => x"ffa5000fffc30000",
    1925 => x"ffa00019ffc30000",
    1926 => x"ffa00019ffc30000",
    1927 => x"ff9b0014ffbd0000",
    1928 => x"00650014ffbd0000",
    1929 => x"006b001bffba0000",
    1930 => x"ff95001bffba0000",
    1931 => x"ff9b0014ffbd0000",
    1932 => x"0062001dffd60000",
    1933 => x"005b000fffc30000",
    1934 => x"ffa5000fffc30000",
    1935 => x"ff9e001dffd60000",
    1936 => x"0053fff8ffd30000",
    1937 => x"0052fffdffc60000",
    1938 => x"ffaefffdffc60000",
    1939 => x"ffadfff8ffd30000",
    1940 => x"006c0019ffb40000",
    1941 => x"006b001bffba0000",
    1942 => x"00650014ffbd0000",
    1943 => x"00650013ffb70000",
    1944 => x"00650013ffb70000",
    1945 => x"006c0019ffb40000",
    1946 => x"ff940019ffb40000",
    1947 => x"ff9b0013ffb70000",
    1948 => x"ff9b0013ffb70000",
    1949 => x"ff9b0014ffbd0000",
    1950 => x"ff95001bffba0000",
    1951 => x"ff940019ffb40000",
    1952 => x"005f000cffbc0000",
    1953 => x"0060000cffb70000",
    1954 => x"0060000cffb70000",
    1955 => x"00650013ffb70000",
    1956 => x"ff9b0013ffb70000",
    1957 => x"ffa0000cffb70000",
    1958 => x"ffa0000cffb70000",
    1959 => x"ffa1000cffbc0000",
    1960 => x"00560003ffbc0000",
    1961 => x"00570003ffb70000",
    1962 => x"00570003ffb70000",
    1963 => x"0060000cffb70000",
    1964 => x"ffa0000cffb70000",
    1965 => x"ffa90003ffb70000",
    1966 => x"ffa90003ffb70000",
    1967 => x"ffaa0003ffbc0000",
    1968 => x"005d0002ffbc0000",
    1969 => x"005e0001ffb70000",
    1970 => x"005e0001ffb70000",
    1971 => x"00570003ffb70000",
    1972 => x"ffa90003ffb70000",
    1973 => x"ffa20001ffb70000",
    1974 => x"ffa20001ffb70000",
    1975 => x"ffa30002ffbc0000",
    1976 => x"0060fffaffbc0000",
    1977 => x"0061fffaffb70000",
    1978 => x"0061fffaffb70000",
    1979 => x"005e0001ffb70000",
    1980 => x"ffa20001ffb70000",
    1981 => x"ff9ffffaffb70000",
    1982 => x"ff9ffffaffb70000",
    1983 => x"ffa0fffaffbc0000",
    1984 => x"005cfff7ffbc0000",
    1985 => x"005cfff7ffb70000",
    1986 => x"005cfff7ffb70000",
    1987 => x"0061fffaffb70000",
    1988 => x"ff9ffffaffb70000",
    1989 => x"ffa4fff7ffb70000",
    1990 => x"ffa4fff7ffb70000",
    1991 => x"ffa4fff7ffbc0000",
    1992 => x"0064fff6ffc30000",
    1993 => x"0064fff7ffbd0000",
    1994 => x"0064fff7ffbd0000",
    1995 => x"005cfff7ffb70000",
    1996 => x"ffa4fff7ffb70000",
    1997 => x"ff9cfff7ffbd0000",
    1998 => x"ff9cfff7ffbd0000",
    1999 => x"ff9cfff6ffc30000",
    2000 => x"0076001effac0000",
    2001 => x"0074001fffb20000",
    2002 => x"006c0019ffb40000",
    2003 => x"0076001effac0000",
    2004 => x"ff8a001effac0000",
    2005 => x"ff940019ffb40000",
    2006 => x"ff8c001fffb20000",
    2007 => x"ff8a001effac0000",
    2008 => x"0087001fffa40000",
    2009 => x"00850021ffa90000",
    2010 => x"0076001effac0000",
    2011 => x"0087001fffa40000",
    2012 => x"ff79001fffa40000",
    2013 => x"ff8a001effac0000",
    2014 => x"ff7b0021ffa90000",
    2015 => x"ff79001fffa40000",
    2016 => x"008f0014ffa30000",
    2017 => x"008c0015ffa90000",
    2018 => x"0087001fffa40000",
    2019 => x"008f0014ffa30000",
    2020 => x"ff710014ffa30000",
    2021 => x"ff79001fffa40000",
    2022 => x"ff740015ffa90000",
    2023 => x"ff710014ffa30000",
    2024 => x"008a0002ffa40000",
    2025 => x"00870003ffa90000",
    2026 => x"008f0014ffa30000",
    2027 => x"008a0002ffa40000",
    2028 => x"ff760002ffa40000",
    2029 => x"ff710014ffa30000",
    2030 => x"ff790003ffa90000",
    2031 => x"ff760002ffa40000",
    2032 => x"0077fff8ffab0000",
    2033 => x"0076fff8ffb10000",
    2034 => x"008a0002ffa40000",
    2035 => x"0077fff8ffab0000",
    2036 => x"ff89fff8ffab0000",
    2037 => x"ff760002ffa40000",
    2038 => x"ff8afff8ffb10000",
    2039 => x"ff89fff8ffab0000",
    2040 => x"0077fff8ffab0000",
    2041 => x"0064fff7ffbd0000",
    2042 => x"ff9cfff7ffbd0000",
    2043 => x"ff89fff8ffab0000",
    2044 => x"00650005ffb60000",
    2045 => x"005e0001ffb70000",
    2046 => x"0061fffaffb70000",
    2047 => x"006bffffffb50000",
    2048 => x"006bffffffb50000",
    2049 => x"00650005ffb60000",
    2050 => x"ff9b0005ffb60000",
    2051 => x"ff95ffffffb50000",
    2052 => x"ff95ffffffb50000",
    2053 => x"ff9ffffaffb70000",
    2054 => x"ffa20001ffb70000",
    2055 => x"ff9b0005ffb60000",
    2056 => x"006d000cffb30000",
    2057 => x"00650005ffb60000",
    2058 => x"006bffffffb50000",
    2059 => x"00720007ffb10000",
    2060 => x"00720007ffb10000",
    2061 => x"006d000cffb30000",
    2062 => x"ff93000cffb30000",
    2063 => x"ff8e0007ffb10000",
    2064 => x"ff8e0007ffb10000",
    2065 => x"ff95ffffffb50000",
    2066 => x"ff9b0005ffb60000",
    2067 => x"ff93000cffb30000",
    2068 => x"00730013ffb10000",
    2069 => x"006d000cffb30000",
    2070 => x"00720007ffb10000",
    2071 => x"0078000effb00000",
    2072 => x"0078000effb00000",
    2073 => x"00730013ffb10000",
    2074 => x"ff8d0013ffb10000",
    2075 => x"ff88000effb00000",
    2076 => x"ff88000effb00000",
    2077 => x"ff8e0007ffb10000",
    2078 => x"ff93000cffb30000",
    2079 => x"ff8d0013ffb10000",
    2080 => x"007b0017ffaf0000",
    2081 => x"00730013ffb10000",
    2082 => x"0078000effb00000",
    2083 => x"007e0010ffaf0000",
    2084 => x"007e0010ffaf0000",
    2085 => x"007b0017ffaf0000",
    2086 => x"ff850017ffaf0000",
    2087 => x"ff820010ffaf0000",
    2088 => x"ff820010ffaf0000",
    2089 => x"ff88000effb00000",
    2090 => x"ff8d0013ffb10000",
    2091 => x"ff850017ffaf0000",
    2092 => x"007b0017ffaf0000",
    2093 => x"0076001effac0000",
    2094 => x"006c0019ffb40000",
    2095 => x"00730013ffb10000",
    2096 => x"ff8d0013ffb10000",
    2097 => x"ff940019ffb40000",
    2098 => x"ff8a001effac0000",
    2099 => x"ff850017ffaf0000",
    2100 => x"00650013ffb70000",
    2101 => x"006d000cffb30000",
    2102 => x"ff93000cffb30000",
    2103 => x"ff9b0013ffb70000",
    2104 => x"0060000cffb70000",
    2105 => x"00650005ffb60000",
    2106 => x"ff9b0005ffb60000",
    2107 => x"ffa0000cffb70000",
    2108 => x"0064fff7ffbd0000",
    2109 => x"006bffffffb50000",
    2110 => x"ff95ffffffb50000",
    2111 => x"ff9cfff7ffbd0000",
    2112 => x"0077fff8ffab0000",
    2113 => x"00720007ffb10000",
    2114 => x"ff8e0007ffb10000",
    2115 => x"ff89fff8ffab0000",
    2116 => x"008a0002ffa40000",
    2117 => x"0078000effb00000",
    2118 => x"ff88000effb00000",
    2119 => x"ff760002ffa40000",
    2120 => x"008f0014ffa30000",
    2121 => x"007e0010ffaf0000",
    2122 => x"ff820010ffaf0000",
    2123 => x"ff710014ffa30000",
    2124 => x"0087001fffa40000",
    2125 => x"007b0017ffaf0000",
    2126 => x"ff850017ffaf0000",
    2127 => x"ff79001fffa40000",
    2128 => x"0076ffefffa30000",
    2129 => x"0076ffedffb60000",
    2130 => x"0058ffe8ffcd0000",
    2131 => x"005affeaffb60000",
    2132 => x"005affeaffb60000",
    2133 => x"0076ffefffa30000",
    2134 => x"ff8affefffa30000",
    2135 => x"ffa6ffeaffb60000",
    2136 => x"ffa6ffeaffb60000",
    2137 => x"ffa8ffe8ffcd0000",
    2138 => x"ff8affedffb60000",
    2139 => x"ff8affefffa30000",
    2140 => x"0095ffffff9f0000",
    2141 => x"0092ffffffaa0000",
    2142 => x"0076ffefffa30000",
    2143 => x"0095ffffff9f0000",
    2144 => x"ff6bffffff9f0000",
    2145 => x"ff8affefffa30000",
    2146 => x"ff6effffffaa0000",
    2147 => x"ff6bffffff9f0000",
    2148 => x"009b001affa20000",
    2149 => x"009a001dffab0000",
    2150 => x"0095ffffff9f0000",
    2151 => x"009b001affa20000",
    2152 => x"ff65001affa20000",
    2153 => x"ff6bffffff9f0000",
    2154 => x"ff66001dffab0000",
    2155 => x"ff65001affa20000",
    2156 => x"008e002eff9d0000",
    2157 => x"008c0032ffab0000",
    2158 => x"009b001affa20000",
    2159 => x"008e002eff9d0000",
    2160 => x"ff72002eff9d0000",
    2161 => x"ff65001affa20000",
    2162 => x"ff740032ffab0000",
    2163 => x"ff72002eff9d0000",
    2164 => x"0074002affa40000",
    2165 => x"0074002fffb80000",
    2166 => x"008e002eff9d0000",
    2167 => x"0074002affa40000",
    2168 => x"ff8c002affa40000",
    2169 => x"ff72002eff9d0000",
    2170 => x"ff8c002fffb80000",
    2171 => x"ff8c002affa40000",
    2172 => x"00620024ffb00000",
    2173 => x"00650027ffc10000",
    2174 => x"0074002affa40000",
    2175 => x"00620024ffb00000",
    2176 => x"ff9e0024ffb00000",
    2177 => x"ff8c002affa40000",
    2178 => x"ff9b0027ffc10000",
    2179 => x"ff9e0024ffb00000",
    2180 => x"0074002affa40000",
    2181 => x"0076ffefffa30000",
    2182 => x"005affeaffb60000",
    2183 => x"00620024ffb00000",
    2184 => x"ff9e0024ffb00000",
    2185 => x"ffa6ffeaffb60000",
    2186 => x"ff8affefffa30000",
    2187 => x"ff8c002affa40000",
    2188 => x"008e002eff9d0000",
    2189 => x"0095ffffff9f0000",
    2190 => x"ff6bffffff9f0000",
    2191 => x"ff72002eff9d0000",
    2192 => x"00620024ffb00000",
    2193 => x"00580017ffa90000",
    2194 => x"ffa80017ffa90000",
    2195 => x"ff9e0024ffb00000",
    2196 => x"005affeaffb60000",
    2197 => x"0049fff7ffaa0000",
    2198 => x"ffb7fff7ffaa0000",
    2199 => x"ffa6ffeaffb60000",
    2200 => x"ffffffffffffffff",
    2201 => x"ffffffffffffffff",

        others => (others => '0'));

begin

PROCESS(clk)
BEGIN
  if (rising_edge(clk)) then
    -- synkron skrivning/läsning port 1
    read_data <= ram(to_integer(read_addr));
  end if;
END PROCESS;

end Behavioral;
